module sample_rom (
	input 		     clk	,
	input 			 ce		,
	input      [5:0] sample	,
	input 	   [7:0] prog	,
	output reg [7:0] d
);

reg [7:0] sample_rom [255:0][63:0];
   
   	//initial
	//	$readmemh("sample_rom.mem", sample_rom );

always @(posedge clk)
	if (ce)
    	d <= sample_rom[prog][sample];

initial begin
	sample_rom[0][0] = 8'd131;
	sample_rom[0][1] = 8'd162;
	sample_rom[0][2] = 8'd188;
	sample_rom[0][3] = 8'd205;
	sample_rom[0][4] = 8'd211;
	sample_rom[0][5] = 8'd208;
	sample_rom[0][6] = 8'd196;
	sample_rom[0][7] = 8'd181;
	sample_rom[0][8] = 8'd164;
	sample_rom[0][9] = 8'd150;
	sample_rom[0][10] = 8'd141;
	sample_rom[0][11] = 8'd134;
	sample_rom[0][12] = 8'd132;
	sample_rom[0][13] = 8'd126;
	sample_rom[0][14] = 8'd119;
	sample_rom[0][15] = 8'd108;
	sample_rom[0][16] = 8'd96;
	sample_rom[0][17] = 8'd82;
	sample_rom[0][18] = 8'd70;
	sample_rom[0][19] = 8'd65;
	sample_rom[0][20] = 8'd68;
	sample_rom[0][21] = 8'd81;
	sample_rom[0][22] = 8'd101;
	sample_rom[0][23] = 8'd125;
	sample_rom[0][24] = 8'd149;
	sample_rom[0][25] = 8'd167;
	sample_rom[0][26] = 8'd178;
	sample_rom[0][27] = 8'd178;
	sample_rom[0][28] = 8'd169;
	sample_rom[0][29] = 8'd154;
	sample_rom[0][30] = 8'd134;
	sample_rom[0][31] = 8'd115;
	sample_rom[0][32] = 8'd103;
	sample_rom[0][33] = 8'd97;
	sample_rom[0][34] = 8'd98;
	sample_rom[0][35] = 8'd105;
	sample_rom[0][36] = 8'd114;
	sample_rom[0][37] = 8'd122;
	sample_rom[0][38] = 8'd127;
	sample_rom[0][39] = 8'd129;
	sample_rom[0][40] = 8'd127;
	sample_rom[0][41] = 8'd126;
	sample_rom[0][42] = 8'd125;
	sample_rom[0][43] = 8'd130;
	sample_rom[0][44] = 8'd142;
	sample_rom[0][45] = 8'd156;
	sample_rom[0][46] = 8'd171;
	sample_rom[0][47] = 8'd186;
	sample_rom[0][48] = 8'd194;
	sample_rom[0][49] = 8'd193;
	sample_rom[0][50] = 8'd182;
	sample_rom[0][51] = 8'd161;
	sample_rom[0][52] = 8'd132;
	sample_rom[0][53] = 8'd102;
	sample_rom[0][54] = 8'd75;
	sample_rom[0][55] = 8'd54;
	sample_rom[0][56] = 8'd45;
	sample_rom[0][57] = 8'd47;
	sample_rom[0][58] = 8'd55;
	sample_rom[0][59] = 8'd71;
	sample_rom[0][60] = 8'd87;
	sample_rom[0][61] = 8'd103;
	sample_rom[0][62] = 8'd114;
	sample_rom[0][63] = 8'd124;
	sample_rom[1][0] = 8'd129;
	sample_rom[1][1] = 8'd167;
	sample_rom[1][2] = 8'd196;
	sample_rom[1][3] = 8'd213;
	sample_rom[1][4] = 8'd219;
	sample_rom[1][5] = 8'd215;
	sample_rom[1][6] = 8'd201;
	sample_rom[1][7] = 8'd185;
	sample_rom[1][8] = 8'd169;
	sample_rom[1][9] = 8'd156;
	sample_rom[1][10] = 8'd147;
	sample_rom[1][11] = 8'd142;
	sample_rom[1][12] = 8'd139;
	sample_rom[1][13] = 8'd135;
	sample_rom[1][14] = 8'd130;
	sample_rom[1][15] = 8'd124;
	sample_rom[1][16] = 8'd118;
	sample_rom[1][17] = 8'd115;
	sample_rom[1][18] = 8'd115;
	sample_rom[1][19] = 8'd120;
	sample_rom[1][20] = 8'd128;
	sample_rom[1][21] = 8'd140;
	sample_rom[1][22] = 8'd150;
	sample_rom[1][23] = 8'd156;
	sample_rom[1][24] = 8'd161;
	sample_rom[1][25] = 8'd160;
	sample_rom[1][26] = 8'd155;
	sample_rom[1][27] = 8'd149;
	sample_rom[1][28] = 8'd140;
	sample_rom[1][29] = 8'd134;
	sample_rom[1][30] = 8'd127;
	sample_rom[1][31] = 8'd124;
	sample_rom[1][32] = 8'd121;
	sample_rom[1][33] = 8'd119;
	sample_rom[1][34] = 8'd119;
	sample_rom[1][35] = 8'd119;
	sample_rom[1][36] = 8'd119;
	sample_rom[1][37] = 8'd117;
	sample_rom[1][38] = 8'd117;
	sample_rom[1][39] = 8'd115;
	sample_rom[1][40] = 8'd113;
	sample_rom[1][41] = 8'd108;
	sample_rom[1][42] = 8'd104;
	sample_rom[1][43] = 8'd103;
	sample_rom[1][44] = 8'd103;
	sample_rom[1][45] = 8'd111;
	sample_rom[1][46] = 8'd121;
	sample_rom[1][47] = 8'd134;
	sample_rom[1][48] = 8'd148;
	sample_rom[1][49] = 8'd159;
	sample_rom[1][50] = 8'd161;
	sample_rom[1][51] = 8'd152;
	sample_rom[1][52] = 8'd136;
	sample_rom[1][53] = 8'd112;
	sample_rom[1][54] = 8'd88;
	sample_rom[1][55] = 8'd63;
	sample_rom[1][56] = 8'd47;
	sample_rom[1][57] = 8'd41;
	sample_rom[1][58] = 8'd43;
	sample_rom[1][59] = 8'd56;
	sample_rom[1][60] = 8'd71;
	sample_rom[1][61] = 8'd88;
	sample_rom[1][62] = 8'd103;
	sample_rom[1][63] = 8'd118;
	sample_rom[2][0] = 8'd130;
	sample_rom[2][1] = 8'd164;
	sample_rom[2][2] = 8'd192;
	sample_rom[2][3] = 8'd214;
	sample_rom[2][4] = 8'd225;
	sample_rom[2][5] = 8'd227;
	sample_rom[2][6] = 8'd223;
	sample_rom[2][7] = 8'd210;
	sample_rom[2][8] = 8'd194;
	sample_rom[2][9] = 8'd178;
	sample_rom[2][10] = 8'd162;
	sample_rom[2][11] = 8'd150;
	sample_rom[2][12] = 8'd141;
	sample_rom[2][13] = 8'd136;
	sample_rom[2][14] = 8'd134;
	sample_rom[2][15] = 8'd133;
	sample_rom[2][16] = 8'd134;
	sample_rom[2][17] = 8'd133;
	sample_rom[2][18] = 8'd138;
	sample_rom[2][19] = 8'd142;
	sample_rom[2][20] = 8'd146;
	sample_rom[2][21] = 8'd151;
	sample_rom[2][22] = 8'd157;
	sample_rom[2][23] = 8'd161;
	sample_rom[2][24] = 8'd163;
	sample_rom[2][25] = 8'd163;
	sample_rom[2][26] = 8'd160;
	sample_rom[2][27] = 8'd154;
	sample_rom[2][28] = 8'd145;
	sample_rom[2][29] = 8'd139;
	sample_rom[2][30] = 8'd133;
	sample_rom[2][31] = 8'd128;
	sample_rom[2][32] = 8'd126;
	sample_rom[2][33] = 8'd128;
	sample_rom[2][34] = 8'd130;
	sample_rom[2][35] = 8'd135;
	sample_rom[2][36] = 8'd136;
	sample_rom[2][37] = 8'd134;
	sample_rom[2][38] = 8'd130;
	sample_rom[2][39] = 8'd123;
	sample_rom[2][40] = 8'd116;
	sample_rom[2][41] = 8'd109;
	sample_rom[2][42] = 8'd102;
	sample_rom[2][43] = 8'd102;
	sample_rom[2][44] = 8'd106;
	sample_rom[2][45] = 8'd116;
	sample_rom[2][46] = 8'd127;
	sample_rom[2][47] = 8'd138;
	sample_rom[2][48] = 8'd149;
	sample_rom[2][49] = 8'd152;
	sample_rom[2][50] = 8'd151;
	sample_rom[2][51] = 8'd141;
	sample_rom[2][52] = 8'd128;
	sample_rom[2][53] = 8'd106;
	sample_rom[2][54] = 8'd86;
	sample_rom[2][55] = 8'd66;
	sample_rom[2][56] = 8'd50;
	sample_rom[2][57] = 8'd42;
	sample_rom[2][58] = 8'd38;
	sample_rom[2][59] = 8'd43;
	sample_rom[2][60] = 8'd53;
	sample_rom[2][61] = 8'd69;
	sample_rom[2][62] = 8'd88;
	sample_rom[2][63] = 8'd108;
	sample_rom[3][0] = 8'd132;
	sample_rom[3][1] = 8'd211;
	sample_rom[3][2] = 8'd241;
	sample_rom[3][3] = 8'd223;
	sample_rom[3][4] = 8'd198;
	sample_rom[3][5] = 8'd191;
	sample_rom[3][6] = 8'd192;
	sample_rom[3][7] = 8'd200;
	sample_rom[3][8] = 8'd215;
	sample_rom[3][9] = 8'd223;
	sample_rom[3][10] = 8'd214;
	sample_rom[3][11] = 8'd191;
	sample_rom[3][12] = 8'd183;
	sample_rom[3][13] = 8'd183;
	sample_rom[3][14] = 8'd184;
	sample_rom[3][15] = 8'd173;
	sample_rom[3][16] = 8'd160;
	sample_rom[3][17] = 8'd143;
	sample_rom[3][18] = 8'd131;
	sample_rom[3][19] = 8'd122;
	sample_rom[3][20] = 8'd130;
	sample_rom[3][21] = 8'd148;
	sample_rom[3][22] = 8'd154;
	sample_rom[3][23] = 8'd145;
	sample_rom[3][24] = 8'd131;
	sample_rom[3][25] = 8'd119;
	sample_rom[3][26] = 8'd119;
	sample_rom[3][27] = 8'd130;
	sample_rom[3][28] = 8'd150;
	sample_rom[3][29] = 8'd163;
	sample_rom[3][30] = 8'd168;
	sample_rom[3][31] = 8'd170;
	sample_rom[3][32] = 8'd176;
	sample_rom[3][33] = 8'd181;
	sample_rom[3][34] = 8'd180;
	sample_rom[3][35] = 8'd171;
	sample_rom[3][36] = 8'd164;
	sample_rom[3][37] = 8'd163;
	sample_rom[3][38] = 8'd165;
	sample_rom[3][39] = 8'd164;
	sample_rom[3][40] = 8'd164;
	sample_rom[3][41] = 8'd167;
	sample_rom[3][42] = 8'd160;
	sample_rom[3][43] = 8'd165;
	sample_rom[3][44] = 8'd167;
	sample_rom[3][45] = 8'd167;
	sample_rom[3][46] = 8'd169;
	sample_rom[3][47] = 8'd164;
	sample_rom[3][48] = 8'd164;
	sample_rom[3][49] = 8'd168;
	sample_rom[3][50] = 8'd164;
	sample_rom[3][51] = 8'd162;
	sample_rom[3][52] = 8'd160;
	sample_rom[3][53] = 8'd160;
	sample_rom[3][54] = 8'd153;
	sample_rom[3][55] = 8'd143;
	sample_rom[3][56] = 8'd149;
	sample_rom[3][57] = 8'd150;
	sample_rom[3][58] = 8'd141;
	sample_rom[3][59] = 8'd135;
	sample_rom[3][60] = 8'd132;
	sample_rom[3][61] = 8'd130;
	sample_rom[3][62] = 8'd128;
	sample_rom[3][63] = 8'd128;
	sample_rom[4][0] = 8'd128;
	sample_rom[4][1] = 8'd128;
	sample_rom[4][2] = 8'd128;
	sample_rom[4][3] = 8'd128;
	sample_rom[4][4] = 8'd128;
	sample_rom[4][5] = 8'd128;
	sample_rom[4][6] = 8'd128;
	sample_rom[4][7] = 8'd128;
	sample_rom[4][8] = 8'd128;
	sample_rom[4][9] = 8'd128;
	sample_rom[4][10] = 8'd128;
	sample_rom[4][11] = 8'd128;
	sample_rom[4][12] = 8'd128;
	sample_rom[4][13] = 8'd128;
	sample_rom[4][14] = 8'd128;
	sample_rom[4][15] = 8'd128;
	sample_rom[4][16] = 8'd128;
	sample_rom[4][17] = 8'd128;
	sample_rom[4][18] = 8'd128;
	sample_rom[4][19] = 8'd128;
	sample_rom[4][20] = 8'd128;
	sample_rom[4][21] = 8'd128;
	sample_rom[4][22] = 8'd128;
	sample_rom[4][23] = 8'd128;
	sample_rom[4][24] = 8'd128;
	sample_rom[4][25] = 8'd128;
	sample_rom[4][26] = 8'd128;
	sample_rom[4][27] = 8'd128;
	sample_rom[4][28] = 8'd128;
	sample_rom[4][29] = 8'd128;
	sample_rom[4][30] = 8'd128;
	sample_rom[4][31] = 8'd128;
	sample_rom[4][32] = 8'd128;
	sample_rom[4][33] = 8'd128;
	sample_rom[4][34] = 8'd128;
	sample_rom[4][35] = 8'd128;
	sample_rom[4][36] = 8'd128;
	sample_rom[4][37] = 8'd128;
	sample_rom[4][38] = 8'd128;
	sample_rom[4][39] = 8'd128;
	sample_rom[4][40] = 8'd128;
	sample_rom[4][41] = 8'd128;
	sample_rom[4][42] = 8'd128;
	sample_rom[4][43] = 8'd128;
	sample_rom[4][44] = 8'd128;
	sample_rom[4][45] = 8'd128;
	sample_rom[4][46] = 8'd128;
	sample_rom[4][47] = 8'd128;
	sample_rom[4][48] = 8'd128;
	sample_rom[4][49] = 8'd128;
	sample_rom[4][50] = 8'd128;
	sample_rom[4][51] = 8'd128;
	sample_rom[4][52] = 8'd128;
	sample_rom[4][53] = 8'd128;
	sample_rom[4][54] = 8'd128;
	sample_rom[4][55] = 8'd128;
	sample_rom[4][56] = 8'd128;
	sample_rom[4][57] = 8'd128;
	sample_rom[4][58] = 8'd128;
	sample_rom[4][59] = 8'd128;
	sample_rom[4][60] = 8'd128;
	sample_rom[4][61] = 8'd128;
	sample_rom[4][62] = 8'd128;
	sample_rom[4][63] = 8'd128;
	sample_rom[5][0] = 8'd130;
	sample_rom[5][1] = 8'd152;
	sample_rom[5][2] = 8'd169;
	sample_rom[5][3] = 8'd185;
	sample_rom[5][4] = 8'd197;
	sample_rom[5][5] = 8'd205;
	sample_rom[5][6] = 8'd206;
	sample_rom[5][7] = 8'd204;
	sample_rom[5][8] = 8'd196;
	sample_rom[5][9] = 8'd185;
	sample_rom[5][10] = 8'd172;
	sample_rom[5][11] = 8'd159;
	sample_rom[5][12] = 8'd145;
	sample_rom[5][13] = 8'd132;
	sample_rom[5][14] = 8'd124;
	sample_rom[5][15] = 8'd119;
	sample_rom[5][16] = 8'd117;
	sample_rom[5][17] = 8'd121;
	sample_rom[5][18] = 8'd130;
	sample_rom[5][19] = 8'd141;
	sample_rom[5][20] = 8'd157;
	sample_rom[5][21] = 8'd173;
	sample_rom[5][22] = 8'd190;
	sample_rom[5][23] = 8'd206;
	sample_rom[5][24] = 8'd218;
	sample_rom[5][25] = 8'd226;
	sample_rom[5][26] = 8'd230;
	sample_rom[5][27] = 8'd230;
	sample_rom[5][28] = 8'd224;
	sample_rom[5][29] = 8'd214;
	sample_rom[5][30] = 8'd199;
	sample_rom[5][31] = 8'd181;
	sample_rom[5][32] = 8'd164;
	sample_rom[5][33] = 8'd146;
	sample_rom[5][34] = 8'd129;
	sample_rom[5][35] = 8'd115;
	sample_rom[5][36] = 8'd105;
	sample_rom[5][37] = 8'd97;
	sample_rom[5][38] = 8'd98;
	sample_rom[5][39] = 8'd101;
	sample_rom[5][40] = 8'd109;
	sample_rom[5][41] = 8'd121;
	sample_rom[5][42] = 8'd135;
	sample_rom[5][43] = 8'd151;
	sample_rom[5][44] = 8'd163;
	sample_rom[5][45] = 8'd177;
	sample_rom[5][46] = 8'd185;
	sample_rom[5][47] = 8'd191;
	sample_rom[5][48] = 8'd193;
	sample_rom[5][49] = 8'd188;
	sample_rom[5][50] = 8'd179;
	sample_rom[5][51] = 8'd167;
	sample_rom[5][52] = 8'd153;
	sample_rom[5][53] = 8'd134;
	sample_rom[5][54] = 8'd116;
	sample_rom[5][55] = 8'd99;
	sample_rom[5][56] = 8'd88;
	sample_rom[5][57] = 8'd78;
	sample_rom[5][58] = 8'd72;
	sample_rom[5][59] = 8'd72;
	sample_rom[5][60] = 8'd77;
	sample_rom[5][61] = 8'd85;
	sample_rom[5][62] = 8'd97;
	sample_rom[5][63] = 8'd113;
	sample_rom[6][0] = 8'd132;
	sample_rom[6][1] = 8'd160;
	sample_rom[6][2] = 8'd185;
	sample_rom[6][3] = 8'd203;
	sample_rom[6][4] = 8'd211;
	sample_rom[6][5] = 8'd211;
	sample_rom[6][6] = 8'd202;
	sample_rom[6][7] = 8'd190;
	sample_rom[6][8] = 8'd177;
	sample_rom[6][9] = 8'd167;
	sample_rom[6][10] = 8'd161;
	sample_rom[6][11] = 8'd160;
	sample_rom[6][12] = 8'd166;
	sample_rom[6][13] = 8'd172;
	sample_rom[6][14] = 8'd178;
	sample_rom[6][15] = 8'd182;
	sample_rom[6][16] = 8'd182;
	sample_rom[6][17] = 8'd176;
	sample_rom[6][18] = 8'd166;
	sample_rom[6][19] = 8'd155;
	sample_rom[6][20] = 8'd146;
	sample_rom[6][21] = 8'd138;
	sample_rom[6][22] = 8'd136;
	sample_rom[6][23] = 8'd140;
	sample_rom[6][24] = 8'd150;
	sample_rom[6][25] = 8'd162;
	sample_rom[6][26] = 8'd174;
	sample_rom[6][27] = 8'd184;
	sample_rom[6][28] = 8'd186;
	sample_rom[6][29] = 8'd181;
	sample_rom[6][30] = 8'd166;
	sample_rom[6][31] = 8'd149;
	sample_rom[6][32] = 8'd126;
	sample_rom[6][33] = 8'd105;
	sample_rom[6][34] = 8'd89;
	sample_rom[6][35] = 8'd82;
	sample_rom[6][36] = 8'd83;
	sample_rom[6][37] = 8'd91;
	sample_rom[6][38] = 8'd108;
	sample_rom[6][39] = 8'd129;
	sample_rom[6][40] = 8'd150;
	sample_rom[6][41] = 8'd167;
	sample_rom[6][42] = 8'd180;
	sample_rom[6][43] = 8'd188;
	sample_rom[6][44] = 8'd188;
	sample_rom[6][45] = 8'd186;
	sample_rom[6][46] = 8'd182;
	sample_rom[6][47] = 8'd181;
	sample_rom[6][48] = 8'd182;
	sample_rom[6][49] = 8'd185;
	sample_rom[6][50] = 8'd193;
	sample_rom[6][51] = 8'd202;
	sample_rom[6][52] = 8'd207;
	sample_rom[6][53] = 8'd209;
	sample_rom[6][54] = 8'd203;
	sample_rom[6][55] = 8'd192;
	sample_rom[6][56] = 8'd175;
	sample_rom[6][57] = 8'd154;
	sample_rom[6][58] = 8'd132;
	sample_rom[6][59] = 8'd114;
	sample_rom[6][60] = 8'd103;
	sample_rom[6][61] = 8'd97;
	sample_rom[6][62] = 8'd103;
	sample_rom[6][63] = 8'd114;
	sample_rom[7][0] = 8'd131;
	sample_rom[7][1] = 8'd176;
	sample_rom[7][2] = 8'd206;
	sample_rom[7][3] = 8'd210;
	sample_rom[7][4] = 8'd188;
	sample_rom[7][5] = 8'd158;
	sample_rom[7][6] = 8'd129;
	sample_rom[7][7] = 8'd114;
	sample_rom[7][8] = 8'd114;
	sample_rom[7][9] = 8'd122;
	sample_rom[7][10] = 8'd126;
	sample_rom[7][11] = 8'd125;
	sample_rom[7][12] = 8'd112;
	sample_rom[7][13] = 8'd99;
	sample_rom[7][14] = 8'd94;
	sample_rom[7][15] = 8'd98;
	sample_rom[7][16] = 8'd112;
	sample_rom[7][17] = 8'd125;
	sample_rom[7][18] = 8'd135;
	sample_rom[7][19] = 8'd134;
	sample_rom[7][20] = 8'd131;
	sample_rom[7][21] = 8'd129;
	sample_rom[7][22] = 8'd137;
	sample_rom[7][23] = 8'd152;
	sample_rom[7][24] = 8'd166;
	sample_rom[7][25] = 8'd171;
	sample_rom[7][26] = 8'd160;
	sample_rom[7][27] = 8'd132;
	sample_rom[7][28] = 8'd97;
	sample_rom[7][29] = 8'd73;
	sample_rom[7][30] = 8'd70;
	sample_rom[7][31] = 8'd93;
	sample_rom[7][32] = 8'd131;
	sample_rom[7][33] = 8'd166;
	sample_rom[7][34] = 8'd186;
	sample_rom[7][35] = 8'd182;
	sample_rom[7][36] = 8'd157;
	sample_rom[7][37] = 8'd123;
	sample_rom[7][38] = 8'd96;
	sample_rom[7][39] = 8'd85;
	sample_rom[7][40] = 8'd91;
	sample_rom[7][41] = 8'd106;
	sample_rom[7][42] = 8'd120;
	sample_rom[7][43] = 8'd129;
	sample_rom[7][44] = 8'd126;
	sample_rom[7][45] = 8'd123;
	sample_rom[7][46] = 8'd123;
	sample_rom[7][47] = 8'd132;
	sample_rom[7][48] = 8'd147;
	sample_rom[7][49] = 8'd159;
	sample_rom[7][50] = 8'd162;
	sample_rom[7][51] = 8'd156;
	sample_rom[7][52] = 8'd143;
	sample_rom[7][53] = 8'd131;
	sample_rom[7][54] = 8'd129;
	sample_rom[7][55] = 8'd134;
	sample_rom[7][56] = 8'd141;
	sample_rom[7][57] = 8'd140;
	sample_rom[7][58] = 8'd126;
	sample_rom[7][59] = 8'd98;
	sample_rom[7][60] = 8'd66;
	sample_rom[7][61] = 8'd47;
	sample_rom[7][62] = 8'd52;
	sample_rom[7][63] = 8'd83;
	sample_rom[8][0] = 8'd132;
	sample_rom[8][1] = 8'd193;
	sample_rom[8][2] = 8'd233;
	sample_rom[8][3] = 8'd245;
	sample_rom[8][4] = 8'd237;
	sample_rom[8][5] = 8'd223;
	sample_rom[8][6] = 8'd211;
	sample_rom[8][7] = 8'd204;
	sample_rom[8][8] = 8'd201;
	sample_rom[8][9] = 8'd196;
	sample_rom[8][10] = 8'd188;
	sample_rom[8][11] = 8'd183;
	sample_rom[8][12] = 8'd177;
	sample_rom[8][13] = 8'd171;
	sample_rom[8][14] = 8'd170;
	sample_rom[8][15] = 8'd172;
	sample_rom[8][16] = 8'd177;
	sample_rom[8][17] = 8'd180;
	sample_rom[8][18] = 8'd179;
	sample_rom[8][19] = 8'd166;
	sample_rom[8][20] = 8'd157;
	sample_rom[8][21] = 8'd146;
	sample_rom[8][22] = 8'd143;
	sample_rom[8][23] = 8'd147;
	sample_rom[8][24] = 8'd149;
	sample_rom[8][25] = 8'd148;
	sample_rom[8][26] = 8'd141;
	sample_rom[8][27] = 8'd130;
	sample_rom[8][28] = 8'd121;
	sample_rom[8][29] = 8'd121;
	sample_rom[8][30] = 8'd124;
	sample_rom[8][31] = 8'd141;
	sample_rom[8][32] = 8'd162;
	sample_rom[8][33] = 8'd178;
	sample_rom[8][34] = 8'd184;
	sample_rom[8][35] = 8'd178;
	sample_rom[8][36] = 8'd166;
	sample_rom[8][37] = 8'd150;
	sample_rom[8][38] = 8'd141;
	sample_rom[8][39] = 8'd139;
	sample_rom[8][40] = 8'd142;
	sample_rom[8][41] = 8'd145;
	sample_rom[8][42] = 8'd142;
	sample_rom[8][43] = 8'd135;
	sample_rom[8][44] = 8'd125;
	sample_rom[8][45] = 8'd115;
	sample_rom[8][46] = 8'd111;
	sample_rom[8][47] = 8'd112;
	sample_rom[8][48] = 8'd120;
	sample_rom[8][49] = 8'd130;
	sample_rom[8][50] = 8'd141;
	sample_rom[8][51] = 8'd142;
	sample_rom[8][52] = 8'd139;
	sample_rom[8][53] = 8'd134;
	sample_rom[8][54] = 8'd129;
	sample_rom[8][55] = 8'd130;
	sample_rom[8][56] = 8'd124;
	sample_rom[8][57] = 8'd109;
	sample_rom[8][58] = 8'd93;
	sample_rom[8][59] = 8'd74;
	sample_rom[8][60] = 8'd62;
	sample_rom[8][61] = 8'd70;
	sample_rom[8][62] = 8'd84;
	sample_rom[8][63] = 8'd107;
	sample_rom[9][0] = 8'd130;
	sample_rom[9][1] = 8'd158;
	sample_rom[9][2] = 8'd180;
	sample_rom[9][3] = 8'd203;
	sample_rom[9][4] = 8'd219;
	sample_rom[9][5] = 8'd231;
	sample_rom[9][6] = 8'd236;
	sample_rom[9][7] = 8'd240;
	sample_rom[9][8] = 8'd236;
	sample_rom[9][9] = 8'd230;
	sample_rom[9][10] = 8'd222;
	sample_rom[9][11] = 8'd210;
	sample_rom[9][12] = 8'd199;
	sample_rom[9][13] = 8'd185;
	sample_rom[9][14] = 8'd171;
	sample_rom[9][15] = 8'd159;
	sample_rom[9][16] = 8'd150;
	sample_rom[9][17] = 8'd139;
	sample_rom[9][18] = 8'd130;
	sample_rom[9][19] = 8'd123;
	sample_rom[9][20] = 8'd116;
	sample_rom[9][21] = 8'd112;
	sample_rom[9][22] = 8'd108;
	sample_rom[9][23] = 8'd108;
	sample_rom[9][24] = 8'd107;
	sample_rom[9][25] = 8'd108;
	sample_rom[9][26] = 8'd112;
	sample_rom[9][27] = 8'd114;
	sample_rom[9][28] = 8'd117;
	sample_rom[9][29] = 8'd121;
	sample_rom[9][30] = 8'd124;
	sample_rom[9][31] = 8'd126;
	sample_rom[9][32] = 8'd125;
	sample_rom[9][33] = 8'd125;
	sample_rom[9][34] = 8'd123;
	sample_rom[9][35] = 8'd123;
	sample_rom[9][36] = 8'd119;
	sample_rom[9][37] = 8'd116;
	sample_rom[9][38] = 8'd113;
	sample_rom[9][39] = 8'd110;
	sample_rom[9][40] = 8'd112;
	sample_rom[9][41] = 8'd111;
	sample_rom[9][42] = 8'd114;
	sample_rom[9][43] = 8'd117;
	sample_rom[9][44] = 8'd120;
	sample_rom[9][45] = 8'd126;
	sample_rom[9][46] = 8'd133;
	sample_rom[9][47] = 8'd142;
	sample_rom[9][48] = 8'd147;
	sample_rom[9][49] = 8'd156;
	sample_rom[9][50] = 8'd166;
	sample_rom[9][51] = 8'd176;
	sample_rom[9][52] = 8'd188;
	sample_rom[9][53] = 8'd197;
	sample_rom[9][54] = 8'd206;
	sample_rom[9][55] = 8'd211;
	sample_rom[9][56] = 8'd217;
	sample_rom[9][57] = 8'd217;
	sample_rom[9][58] = 8'd218;
	sample_rom[9][59] = 8'd210;
	sample_rom[9][60] = 8'd200;
	sample_rom[9][61] = 8'd185;
	sample_rom[9][62] = 8'd166;
	sample_rom[9][63] = 8'd149;
	sample_rom[10][0] = 8'd130;
	sample_rom[10][1] = 8'd161;
	sample_rom[10][2] = 8'd187;
	sample_rom[10][3] = 8'd209;
	sample_rom[10][4] = 8'd224;
	sample_rom[10][5] = 8'd234;
	sample_rom[10][6] = 8'd241;
	sample_rom[10][7] = 8'd239;
	sample_rom[10][8] = 8'd234;
	sample_rom[10][9] = 8'd225;
	sample_rom[10][10] = 8'd215;
	sample_rom[10][11] = 8'd201;
	sample_rom[10][12] = 8'd186;
	sample_rom[10][13] = 8'd169;
	sample_rom[10][14] = 8'd156;
	sample_rom[10][15] = 8'd139;
	sample_rom[10][16] = 8'd128;
	sample_rom[10][17] = 8'd116;
	sample_rom[10][18] = 8'd112;
	sample_rom[10][19] = 8'd109;
	sample_rom[10][20] = 8'd110;
	sample_rom[10][21] = 8'd112;
	sample_rom[10][22] = 8'd114;
	sample_rom[10][23] = 8'd120;
	sample_rom[10][24] = 8'd124;
	sample_rom[10][25] = 8'd128;
	sample_rom[10][26] = 8'd132;
	sample_rom[10][27] = 8'd138;
	sample_rom[10][28] = 8'd141;
	sample_rom[10][29] = 8'd142;
	sample_rom[10][30] = 8'd141;
	sample_rom[10][31] = 8'd142;
	sample_rom[10][32] = 8'd143;
	sample_rom[10][33] = 8'd140;
	sample_rom[10][34] = 8'd139;
	sample_rom[10][35] = 8'd137;
	sample_rom[10][36] = 8'd137;
	sample_rom[10][37] = 8'd131;
	sample_rom[10][38] = 8'd128;
	sample_rom[10][39] = 8'd124;
	sample_rom[10][40] = 8'd120;
	sample_rom[10][41] = 8'd115;
	sample_rom[10][42] = 8'd112;
	sample_rom[10][43] = 8'd110;
	sample_rom[10][44] = 8'd110;
	sample_rom[10][45] = 8'd110;
	sample_rom[10][46] = 8'd113;
	sample_rom[10][47] = 8'd118;
	sample_rom[10][48] = 8'd123;
	sample_rom[10][49] = 8'd129;
	sample_rom[10][50] = 8'd138;
	sample_rom[10][51] = 8'd147;
	sample_rom[10][52] = 8'd158;
	sample_rom[10][53] = 8'd168;
	sample_rom[10][54] = 8'd179;
	sample_rom[10][55] = 8'd189;
	sample_rom[10][56] = 8'd195;
	sample_rom[10][57] = 8'd198;
	sample_rom[10][58] = 8'd200;
	sample_rom[10][59] = 8'd196;
	sample_rom[10][60] = 8'd185;
	sample_rom[10][61] = 8'd172;
	sample_rom[10][62] = 8'd159;
	sample_rom[10][63] = 8'd143;
	sample_rom[11][0] = 8'd129;
	sample_rom[11][1] = 8'd186;
	sample_rom[11][2] = 8'd223;
	sample_rom[11][3] = 8'd237;
	sample_rom[11][4] = 8'd229;
	sample_rom[11][5] = 8'd210;
	sample_rom[11][6] = 8'd178;
	sample_rom[11][7] = 8'd152;
	sample_rom[11][8] = 8'd123;
	sample_rom[11][9] = 8'd102;
	sample_rom[11][10] = 8'd96;
	sample_rom[11][11] = 8'd98;
	sample_rom[11][12] = 8'd108;
	sample_rom[11][13] = 8'd121;
	sample_rom[11][14] = 8'd130;
	sample_rom[11][15] = 8'd136;
	sample_rom[11][16] = 8'd139;
	sample_rom[11][17] = 8'd140;
	sample_rom[11][18] = 8'd136;
	sample_rom[11][19] = 8'd129;
	sample_rom[11][20] = 8'd124;
	sample_rom[11][21] = 8'd123;
	sample_rom[11][22] = 8'd119;
	sample_rom[11][23] = 8'd122;
	sample_rom[11][24] = 8'd121;
	sample_rom[11][25] = 8'd123;
	sample_rom[11][26] = 8'd124;
	sample_rom[11][27] = 8'd128;
	sample_rom[11][28] = 8'd135;
	sample_rom[11][29] = 8'd138;
	sample_rom[11][30] = 8'd146;
	sample_rom[11][31] = 8'd147;
	sample_rom[11][32] = 8'd148;
	sample_rom[11][33] = 8'd147;
	sample_rom[11][34] = 8'd144;
	sample_rom[11][35] = 8'd142;
	sample_rom[11][36] = 8'd134;
	sample_rom[11][37] = 8'd135;
	sample_rom[11][38] = 8'd128;
	sample_rom[11][39] = 8'd121;
	sample_rom[11][40] = 8'd116;
	sample_rom[11][41] = 8'd113;
	sample_rom[11][42] = 8'd119;
	sample_rom[11][43] = 8'd119;
	sample_rom[11][44] = 8'd127;
	sample_rom[11][45] = 8'd134;
	sample_rom[11][46] = 8'd140;
	sample_rom[11][47] = 8'd140;
	sample_rom[11][48] = 8'd142;
	sample_rom[11][49] = 8'd136;
	sample_rom[11][50] = 8'd125;
	sample_rom[11][51] = 8'd112;
	sample_rom[11][52] = 8'd104;
	sample_rom[11][53] = 8'd93;
	sample_rom[11][54] = 8'd96;
	sample_rom[11][55] = 8'd106;
	sample_rom[11][56] = 8'd128;
	sample_rom[11][57] = 8'd157;
	sample_rom[11][58] = 8'd188;
	sample_rom[11][59] = 8'd207;
	sample_rom[11][60] = 8'd216;
	sample_rom[11][61] = 8'd205;
	sample_rom[11][62] = 8'd180;
	sample_rom[11][63] = 8'd157;
	sample_rom[12][0] = 8'd131;
	sample_rom[12][1] = 8'd160;
	sample_rom[12][2] = 8'd184;
	sample_rom[12][3] = 8'd206;
	sample_rom[12][4] = 8'd223;
	sample_rom[12][5] = 8'd236;
	sample_rom[12][6] = 8'd242;
	sample_rom[12][7] = 8'd244;
	sample_rom[12][8] = 8'd240;
	sample_rom[12][9] = 8'd231;
	sample_rom[12][10] = 8'd220;
	sample_rom[12][11] = 8'd205;
	sample_rom[12][12] = 8'd190;
	sample_rom[12][13] = 8'd172;
	sample_rom[12][14] = 8'd158;
	sample_rom[12][15] = 8'd143;
	sample_rom[12][16] = 8'd133;
	sample_rom[12][17] = 8'd124;
	sample_rom[12][18] = 8'd117;
	sample_rom[12][19] = 8'd114;
	sample_rom[12][20] = 8'd114;
	sample_rom[12][21] = 8'd114;
	sample_rom[12][22] = 8'd115;
	sample_rom[12][23] = 8'd119;
	sample_rom[12][24] = 8'd123;
	sample_rom[12][25] = 8'd125;
	sample_rom[12][26] = 8'd129;
	sample_rom[12][27] = 8'd131;
	sample_rom[12][28] = 8'd134;
	sample_rom[12][29] = 8'd135;
	sample_rom[12][30] = 8'd135;
	sample_rom[12][31] = 8'd136;
	sample_rom[12][32] = 8'd136;
	sample_rom[12][33] = 8'd136;
	sample_rom[12][34] = 8'd135;
	sample_rom[12][35] = 8'd134;
	sample_rom[12][36] = 8'd133;
	sample_rom[12][37] = 8'd131;
	sample_rom[12][38] = 8'd129;
	sample_rom[12][39] = 8'd124;
	sample_rom[12][40] = 8'd123;
	sample_rom[12][41] = 8'd118;
	sample_rom[12][42] = 8'd117;
	sample_rom[12][43] = 8'd114;
	sample_rom[12][44] = 8'd114;
	sample_rom[12][45] = 8'd115;
	sample_rom[12][46] = 8'd120;
	sample_rom[12][47] = 8'd126;
	sample_rom[12][48] = 8'd134;
	sample_rom[12][49] = 8'd146;
	sample_rom[12][50] = 8'd160;
	sample_rom[12][51] = 8'd175;
	sample_rom[12][52] = 8'd192;
	sample_rom[12][53] = 8'd207;
	sample_rom[12][54] = 8'd221;
	sample_rom[12][55] = 8'd232;
	sample_rom[12][56] = 8'd239;
	sample_rom[12][57] = 8'd242;
	sample_rom[12][58] = 8'd240;
	sample_rom[12][59] = 8'd231;
	sample_rom[12][60] = 8'd219;
	sample_rom[12][61] = 8'd199;
	sample_rom[12][62] = 8'd177;
	sample_rom[12][63] = 8'd153;
	sample_rom[13][0] = 8'd134;
	sample_rom[13][1] = 8'd162;
	sample_rom[13][2] = 8'd157;
	sample_rom[13][3] = 8'd229;
	sample_rom[13][4] = 8'd132;
	sample_rom[13][5] = 8'd165;
	sample_rom[13][6] = 8'd165;
	sample_rom[13][7] = 8'd87;
	sample_rom[13][8] = 8'd71;
	sample_rom[13][9] = 8'd167;
	sample_rom[13][10] = 8'd240;
	sample_rom[13][11] = 8'd200;
	sample_rom[13][12] = 8'd135;
	sample_rom[13][13] = 8'd148;
	sample_rom[13][14] = 8'd201;
	sample_rom[13][15] = 8'd208;
	sample_rom[13][16] = 8'd175;
	sample_rom[13][17] = 8'd148;
	sample_rom[13][18] = 8'd127;
	sample_rom[13][19] = 8'd87;
	sample_rom[13][20] = 8'd60;
	sample_rom[13][21] = 8'd82;
	sample_rom[13][22] = 8'd138;
	sample_rom[13][23] = 8'd166;
	sample_rom[13][24] = 8'd158;
	sample_rom[13][25] = 8'd152;
	sample_rom[13][26] = 8'd147;
	sample_rom[13][27] = 8'd110;
	sample_rom[13][28] = 8'd51;
	sample_rom[13][29] = 8'd30;
	sample_rom[13][30] = 8'd76;
	sample_rom[13][31] = 8'd141;
	sample_rom[13][32] = 8'd156;
	sample_rom[13][33] = 8'd128;
	sample_rom[13][34] = 8'd119;
	sample_rom[13][35] = 8'd157;
	sample_rom[13][36] = 8'd170;
	sample_rom[13][37] = 8'd141;
	sample_rom[13][38] = 8'd108;
	sample_rom[13][39] = 8'd121;
	sample_rom[13][40] = 8'd152;
	sample_rom[13][41] = 8'd152;
	sample_rom[13][42] = 8'd114;
	sample_rom[13][43] = 8'd91;
	sample_rom[13][44] = 8'd117;
	sample_rom[13][45] = 8'd163;
	sample_rom[13][46] = 8'd188;
	sample_rom[13][47] = 8'd171;
	sample_rom[13][48] = 8'd135;
	sample_rom[13][49] = 8'd97;
	sample_rom[13][50] = 8'd88;
	sample_rom[13][51] = 8'd103;
	sample_rom[13][52] = 8'd122;
	sample_rom[13][53] = 8'd128;
	sample_rom[13][54] = 8'd144;
	sample_rom[13][55] = 8'd157;
	sample_rom[13][56] = 8'd150;
	sample_rom[13][57] = 8'd102;
	sample_rom[13][58] = 8'd68;
	sample_rom[13][59] = 8'd90;
	sample_rom[13][60] = 8'd133;
	sample_rom[13][61] = 8'd121;
	sample_rom[13][62] = 8'd59;
	sample_rom[13][63] = 8'd49;
	sample_rom[14][0] = 8'd132;
	sample_rom[14][1] = 8'd180;
	sample_rom[14][2] = 8'd217;
	sample_rom[14][3] = 8'd242;
	sample_rom[14][4] = 8'd251;
	sample_rom[14][5] = 8'd253;
	sample_rom[14][6] = 8'd250;
	sample_rom[14][7] = 8'd239;
	sample_rom[14][8] = 8'd224;
	sample_rom[14][9] = 8'd209;
	sample_rom[14][10] = 8'd201;
	sample_rom[14][11] = 8'd194;
	sample_rom[14][12] = 8'd195;
	sample_rom[14][13] = 8'd189;
	sample_rom[14][14] = 8'd187;
	sample_rom[14][15] = 8'd182;
	sample_rom[14][16] = 8'd178;
	sample_rom[14][17] = 8'd170;
	sample_rom[14][18] = 8'd168;
	sample_rom[14][19] = 8'd161;
	sample_rom[14][20] = 8'd158;
	sample_rom[14][21] = 8'd153;
	sample_rom[14][22] = 8'd152;
	sample_rom[14][23] = 8'd153;
	sample_rom[14][24] = 8'd152;
	sample_rom[14][25] = 8'd148;
	sample_rom[14][26] = 8'd135;
	sample_rom[14][27] = 8'd127;
	sample_rom[14][28] = 8'd113;
	sample_rom[14][29] = 8'd105;
	sample_rom[14][30] = 8'd99;
	sample_rom[14][31] = 8'd97;
	sample_rom[14][32] = 8'd100;
	sample_rom[14][33] = 8'd106;
	sample_rom[14][34] = 8'd114;
	sample_rom[14][35] = 8'd122;
	sample_rom[14][36] = 8'd131;
	sample_rom[14][37] = 8'd135;
	sample_rom[14][38] = 8'd141;
	sample_rom[14][39] = 8'd144;
	sample_rom[14][40] = 8'd144;
	sample_rom[14][41] = 8'd142;
	sample_rom[14][42] = 8'd142;
	sample_rom[14][43] = 8'd141;
	sample_rom[14][44] = 8'd145;
	sample_rom[14][45] = 8'd148;
	sample_rom[14][46] = 8'd143;
	sample_rom[14][47] = 8'd134;
	sample_rom[14][48] = 8'd125;
	sample_rom[14][49] = 8'd117;
	sample_rom[14][50] = 8'd111;
	sample_rom[14][51] = 8'd109;
	sample_rom[14][52] = 8'd107;
	sample_rom[14][53] = 8'd104;
	sample_rom[14][54] = 8'd106;
	sample_rom[14][55] = 8'd111;
	sample_rom[14][56] = 8'd118;
	sample_rom[14][57] = 8'd122;
	sample_rom[14][58] = 8'd125;
	sample_rom[14][59] = 8'd128;
	sample_rom[14][60] = 8'd129;
	sample_rom[14][61] = 8'd134;
	sample_rom[14][62] = 8'd136;
	sample_rom[14][63] = 8'd133;
	sample_rom[15][0] = 8'd131;
	sample_rom[15][1] = 8'd164;
	sample_rom[15][2] = 8'd191;
	sample_rom[15][3] = 8'd216;
	sample_rom[15][4] = 8'd233;
	sample_rom[15][5] = 8'd243;
	sample_rom[15][6] = 8'd246;
	sample_rom[15][7] = 8'd239;
	sample_rom[15][8] = 8'd231;
	sample_rom[15][9] = 8'd214;
	sample_rom[15][10] = 8'd194;
	sample_rom[15][11] = 8'd174;
	sample_rom[15][12] = 8'd154;
	sample_rom[15][13] = 8'd129;
	sample_rom[15][14] = 8'd110;
	sample_rom[15][15] = 8'd95;
	sample_rom[15][16] = 8'd83;
	sample_rom[15][17] = 8'd73;
	sample_rom[15][18] = 8'd73;
	sample_rom[15][19] = 8'd74;
	sample_rom[15][20] = 8'd83;
	sample_rom[15][21] = 8'd93;
	sample_rom[15][22] = 8'd107;
	sample_rom[15][23] = 8'd121;
	sample_rom[15][24] = 8'd138;
	sample_rom[15][25] = 8'd153;
	sample_rom[15][26] = 8'd163;
	sample_rom[15][27] = 8'd174;
	sample_rom[15][28] = 8'd184;
	sample_rom[15][29] = 8'd187;
	sample_rom[15][30] = 8'd188;
	sample_rom[15][31] = 8'd189;
	sample_rom[15][32] = 8'd185;
	sample_rom[15][33] = 8'd178;
	sample_rom[15][34] = 8'd169;
	sample_rom[15][35] = 8'd160;
	sample_rom[15][36] = 8'd152;
	sample_rom[15][37] = 8'd141;
	sample_rom[15][38] = 8'd134;
	sample_rom[15][39] = 8'd127;
	sample_rom[15][40] = 8'd122;
	sample_rom[15][41] = 8'd119;
	sample_rom[15][42] = 8'd117;
	sample_rom[15][43] = 8'd118;
	sample_rom[15][44] = 8'd119;
	sample_rom[15][45] = 8'd122;
	sample_rom[15][46] = 8'd125;
	sample_rom[15][47] = 8'd132;
	sample_rom[15][48] = 8'd137;
	sample_rom[15][49] = 8'd140;
	sample_rom[15][50] = 8'd144;
	sample_rom[15][51] = 8'd146;
	sample_rom[15][52] = 8'd147;
	sample_rom[15][53] = 8'd145;
	sample_rom[15][54] = 8'd144;
	sample_rom[15][55] = 8'd140;
	sample_rom[15][56] = 8'd139;
	sample_rom[15][57] = 8'd137;
	sample_rom[15][58] = 8'd135;
	sample_rom[15][59] = 8'd136;
	sample_rom[15][60] = 8'd134;
	sample_rom[15][61] = 8'd134;
	sample_rom[15][62] = 8'd132;
	sample_rom[15][63] = 8'd132;
	sample_rom[16][0] = 8'd128;
	sample_rom[16][1] = 8'd190;
	sample_rom[16][2] = 8'd222;
	sample_rom[16][3] = 8'd222;
	sample_rom[16][4] = 8'd203;
	sample_rom[16][5] = 8'd180;
	sample_rom[16][6] = 8'd162;
	sample_rom[16][7] = 8'd146;
	sample_rom[16][8] = 8'd142;
	sample_rom[16][9] = 8'd146;
	sample_rom[16][10] = 8'd149;
	sample_rom[16][11] = 8'd148;
	sample_rom[16][12] = 8'd143;
	sample_rom[16][13] = 8'd132;
	sample_rom[16][14] = 8'd128;
	sample_rom[16][15] = 8'd131;
	sample_rom[16][16] = 8'd135;
	sample_rom[16][17] = 8'd144;
	sample_rom[16][18] = 8'd154;
	sample_rom[16][19] = 8'd158;
	sample_rom[16][20] = 8'd157;
	sample_rom[16][21] = 8'd150;
	sample_rom[16][22] = 8'd146;
	sample_rom[16][23] = 8'd134;
	sample_rom[16][24] = 8'd127;
	sample_rom[16][25] = 8'd123;
	sample_rom[16][26] = 8'd123;
	sample_rom[16][27] = 8'd128;
	sample_rom[16][28] = 8'd131;
	sample_rom[16][29] = 8'd132;
	sample_rom[16][30] = 8'd137;
	sample_rom[16][31] = 8'd136;
	sample_rom[16][32] = 8'd135;
	sample_rom[16][33] = 8'd141;
	sample_rom[16][34] = 8'd147;
	sample_rom[16][35] = 8'd146;
	sample_rom[16][36] = 8'd146;
	sample_rom[16][37] = 8'd144;
	sample_rom[16][38] = 8'd151;
	sample_rom[16][39] = 8'd147;
	sample_rom[16][40] = 8'd146;
	sample_rom[16][41] = 8'd138;
	sample_rom[16][42] = 8'd135;
	sample_rom[16][43] = 8'd131;
	sample_rom[16][44] = 8'd137;
	sample_rom[16][45] = 8'd136;
	sample_rom[16][46] = 8'd129;
	sample_rom[16][47] = 8'd128;
	sample_rom[16][48] = 8'd125;
	sample_rom[16][49] = 8'd119;
	sample_rom[16][50] = 8'd117;
	sample_rom[16][51] = 8'd114;
	sample_rom[16][52] = 8'd118;
	sample_rom[16][53] = 8'd123;
	sample_rom[16][54] = 8'd131;
	sample_rom[16][55] = 8'd134;
	sample_rom[16][56] = 8'd138;
	sample_rom[16][57] = 8'd137;
	sample_rom[16][58] = 8'd131;
	sample_rom[16][59] = 8'd127;
	sample_rom[16][60] = 8'd125;
	sample_rom[16][61] = 8'd130;
	sample_rom[16][62] = 8'd130;
	sample_rom[16][63] = 8'd128;
	sample_rom[17][0] = 8'd131;
	sample_rom[17][1] = 8'd145;
	sample_rom[17][2] = 8'd157;
	sample_rom[17][3] = 8'd168;
	sample_rom[17][4] = 8'd179;
	sample_rom[17][5] = 8'd190;
	sample_rom[17][6] = 8'd200;
	sample_rom[17][7] = 8'd209;
	sample_rom[17][8] = 8'd216;
	sample_rom[17][9] = 8'd223;
	sample_rom[17][10] = 8'd228;
	sample_rom[17][11] = 8'd232;
	sample_rom[17][12] = 8'd235;
	sample_rom[17][13] = 8'd236;
	sample_rom[17][14] = 8'd237;
	sample_rom[17][15] = 8'd237;
	sample_rom[17][16] = 8'd235;
	sample_rom[17][17] = 8'd231;
	sample_rom[17][18] = 8'd228;
	sample_rom[17][19] = 8'd224;
	sample_rom[17][20] = 8'd219;
	sample_rom[17][21] = 8'd216;
	sample_rom[17][22] = 8'd209;
	sample_rom[17][23] = 8'd203;
	sample_rom[17][24] = 8'd198;
	sample_rom[17][25] = 8'd192;
	sample_rom[17][26] = 8'd186;
	sample_rom[17][27] = 8'd181;
	sample_rom[17][28] = 8'd175;
	sample_rom[17][29] = 8'd169;
	sample_rom[17][30] = 8'd166;
	sample_rom[17][31] = 8'd161;
	sample_rom[17][32] = 8'd158;
	sample_rom[17][33] = 8'd154;
	sample_rom[17][34] = 8'd150;
	sample_rom[17][35] = 8'd148;
	sample_rom[17][36] = 8'd147;
	sample_rom[17][37] = 8'd142;
	sample_rom[17][38] = 8'd141;
	sample_rom[17][39] = 8'd140;
	sample_rom[17][40] = 8'd138;
	sample_rom[17][41] = 8'd137;
	sample_rom[17][42] = 8'd135;
	sample_rom[17][43] = 8'd133;
	sample_rom[17][44] = 8'd132;
	sample_rom[17][45] = 8'd130;
	sample_rom[17][46] = 8'd130;
	sample_rom[17][47] = 8'd128;
	sample_rom[17][48] = 8'd129;
	sample_rom[17][49] = 8'd127;
	sample_rom[17][50] = 8'd126;
	sample_rom[17][51] = 8'd126;
	sample_rom[17][52] = 8'd125;
	sample_rom[17][53] = 8'd125;
	sample_rom[17][54] = 8'd124;
	sample_rom[17][55] = 8'd122;
	sample_rom[17][56] = 8'd122;
	sample_rom[17][57] = 8'd124;
	sample_rom[17][58] = 8'd124;
	sample_rom[17][59] = 8'd125;
	sample_rom[17][60] = 8'd126;
	sample_rom[17][61] = 8'd126;
	sample_rom[17][62] = 8'd125;
	sample_rom[17][63] = 8'd127;
	sample_rom[18][0] = 8'd131;
	sample_rom[18][1] = 8'd150;
	sample_rom[18][2] = 8'd165;
	sample_rom[18][3] = 8'd181;
	sample_rom[18][4] = 8'd195;
	sample_rom[18][5] = 8'd208;
	sample_rom[18][6] = 8'd218;
	sample_rom[18][7] = 8'd226;
	sample_rom[18][8] = 8'd230;
	sample_rom[18][9] = 8'd233;
	sample_rom[18][10] = 8'd235;
	sample_rom[18][11] = 8'd232;
	sample_rom[18][12] = 8'd228;
	sample_rom[18][13] = 8'd222;
	sample_rom[18][14] = 8'd216;
	sample_rom[18][15] = 8'd207;
	sample_rom[18][16] = 8'd196;
	sample_rom[18][17] = 8'd184;
	sample_rom[18][18] = 8'd174;
	sample_rom[18][19] = 8'd162;
	sample_rom[18][20] = 8'd154;
	sample_rom[18][21] = 8'd142;
	sample_rom[18][22] = 8'd134;
	sample_rom[18][23] = 8'd127;
	sample_rom[18][24] = 8'd119;
	sample_rom[18][25] = 8'd114;
	sample_rom[18][26] = 8'd111;
	sample_rom[18][27] = 8'd107;
	sample_rom[18][28] = 8'd105;
	sample_rom[18][29] = 8'd106;
	sample_rom[18][30] = 8'd105;
	sample_rom[18][31] = 8'd107;
	sample_rom[18][32] = 8'd109;
	sample_rom[18][33] = 8'd110;
	sample_rom[18][34] = 8'd113;
	sample_rom[18][35] = 8'd117;
	sample_rom[18][36] = 8'd119;
	sample_rom[18][37] = 8'd120;
	sample_rom[18][38] = 8'd123;
	sample_rom[18][39] = 8'd123;
	sample_rom[18][40] = 8'd126;
	sample_rom[18][41] = 8'd126;
	sample_rom[18][42] = 8'd128;
	sample_rom[18][43] = 8'd128;
	sample_rom[18][44] = 8'd130;
	sample_rom[18][45] = 8'd128;
	sample_rom[18][46] = 8'd130;
	sample_rom[18][47] = 8'd129;
	sample_rom[18][48] = 8'd129;
	sample_rom[18][49] = 8'd128;
	sample_rom[18][50] = 8'd128;
	sample_rom[18][51] = 8'd128;
	sample_rom[18][52] = 8'd129;
	sample_rom[18][53] = 8'd128;
	sample_rom[18][54] = 8'd129;
	sample_rom[18][55] = 8'd129;
	sample_rom[18][56] = 8'd129;
	sample_rom[18][57] = 8'd129;
	sample_rom[18][58] = 8'd129;
	sample_rom[18][59] = 8'd130;
	sample_rom[18][60] = 8'd129;
	sample_rom[18][61] = 8'd129;
	sample_rom[18][62] = 8'd127;
	sample_rom[18][63] = 8'd128;
	sample_rom[19][0] = 8'd129;
	sample_rom[19][1] = 8'd168;
	sample_rom[19][2] = 8'd197;
	sample_rom[19][3] = 8'd225;
	sample_rom[19][4] = 8'd238;
	sample_rom[19][5] = 8'd243;
	sample_rom[19][6] = 8'd237;
	sample_rom[19][7] = 8'd228;
	sample_rom[19][8] = 8'd215;
	sample_rom[19][9] = 8'd197;
	sample_rom[19][10] = 8'd183;
	sample_rom[19][11] = 8'd168;
	sample_rom[19][12] = 8'd155;
	sample_rom[19][13] = 8'd146;
	sample_rom[19][14] = 8'd138;
	sample_rom[19][15] = 8'd132;
	sample_rom[19][16] = 8'd129;
	sample_rom[19][17] = 8'd128;
	sample_rom[19][18] = 8'd129;
	sample_rom[19][19] = 8'd128;
	sample_rom[19][20] = 8'd125;
	sample_rom[19][21] = 8'd127;
	sample_rom[19][22] = 8'd123;
	sample_rom[19][23] = 8'd118;
	sample_rom[19][24] = 8'd116;
	sample_rom[19][25] = 8'd110;
	sample_rom[19][26] = 8'd110;
	sample_rom[19][27] = 8'd109;
	sample_rom[19][28] = 8'd109;
	sample_rom[19][29] = 8'd110;
	sample_rom[19][30] = 8'd114;
	sample_rom[19][31] = 8'd117;
	sample_rom[19][32] = 8'd119;
	sample_rom[19][33] = 8'd121;
	sample_rom[19][34] = 8'd124;
	sample_rom[19][35] = 8'd128;
	sample_rom[19][36] = 8'd126;
	sample_rom[19][37] = 8'd125;
	sample_rom[19][38] = 8'd125;
	sample_rom[19][39] = 8'd124;
	sample_rom[19][40] = 8'd121;
	sample_rom[19][41] = 8'd120;
	sample_rom[19][42] = 8'd119;
	sample_rom[19][43] = 8'd117;
	sample_rom[19][44] = 8'd123;
	sample_rom[19][45] = 8'd126;
	sample_rom[19][46] = 8'd127;
	sample_rom[19][47] = 8'd130;
	sample_rom[19][48] = 8'd134;
	sample_rom[19][49] = 8'd134;
	sample_rom[19][50] = 8'd132;
	sample_rom[19][51] = 8'd132;
	sample_rom[19][52] = 8'd133;
	sample_rom[19][53] = 8'd130;
	sample_rom[19][54] = 8'd132;
	sample_rom[19][55] = 8'd132;
	sample_rom[19][56] = 8'd134;
	sample_rom[19][57] = 8'd135;
	sample_rom[19][58] = 8'd133;
	sample_rom[19][59] = 8'd134;
	sample_rom[19][60] = 8'd129;
	sample_rom[19][61] = 8'd129;
	sample_rom[19][62] = 8'd127;
	sample_rom[19][63] = 8'd127;
	sample_rom[20][0] = 8'd131;
	sample_rom[20][1] = 8'd176;
	sample_rom[20][2] = 8'd211;
	sample_rom[20][3] = 8'd235;
	sample_rom[20][4] = 8'd244;
	sample_rom[20][5] = 8'd243;
	sample_rom[20][6] = 8'd232;
	sample_rom[20][7] = 8'd217;
	sample_rom[20][8] = 8'd199;
	sample_rom[20][9] = 8'd181;
	sample_rom[20][10] = 8'd162;
	sample_rom[20][11] = 8'd151;
	sample_rom[20][12] = 8'd141;
	sample_rom[20][13] = 8'd131;
	sample_rom[20][14] = 8'd128;
	sample_rom[20][15] = 8'd127;
	sample_rom[20][16] = 8'd125;
	sample_rom[20][17] = 8'd124;
	sample_rom[20][18] = 8'd126;
	sample_rom[20][19] = 8'd123;
	sample_rom[20][20] = 8'd122;
	sample_rom[20][21] = 8'd122;
	sample_rom[20][22] = 8'd121;
	sample_rom[20][23] = 8'd122;
	sample_rom[20][24] = 8'd124;
	sample_rom[20][25] = 8'd123;
	sample_rom[20][26] = 8'd118;
	sample_rom[20][27] = 8'd114;
	sample_rom[20][28] = 8'd109;
	sample_rom[20][29] = 8'd111;
	sample_rom[20][30] = 8'd112;
	sample_rom[20][31] = 8'd118;
	sample_rom[20][32] = 8'd123;
	sample_rom[20][33] = 8'd129;
	sample_rom[20][34] = 8'd130;
	sample_rom[20][35] = 8'd129;
	sample_rom[20][36] = 8'd130;
	sample_rom[20][37] = 8'd127;
	sample_rom[20][38] = 8'd124;
	sample_rom[20][39] = 8'd120;
	sample_rom[20][40] = 8'd121;
	sample_rom[20][41] = 8'd120;
	sample_rom[20][42] = 8'd120;
	sample_rom[20][43] = 8'd125;
	sample_rom[20][44] = 8'd128;
	sample_rom[20][45] = 8'd130;
	sample_rom[20][46] = 8'd133;
	sample_rom[20][47] = 8'd132;
	sample_rom[20][48] = 8'd129;
	sample_rom[20][49] = 8'd129;
	sample_rom[20][50] = 8'd128;
	sample_rom[20][51] = 8'd126;
	sample_rom[20][52] = 8'd130;
	sample_rom[20][53] = 8'd129;
	sample_rom[20][54] = 8'd132;
	sample_rom[20][55] = 8'd130;
	sample_rom[20][56] = 8'd133;
	sample_rom[20][57] = 8'd132;
	sample_rom[20][58] = 8'd132;
	sample_rom[20][59] = 8'd133;
	sample_rom[20][60] = 8'd130;
	sample_rom[20][61] = 8'd132;
	sample_rom[20][62] = 8'd130;
	sample_rom[20][63] = 8'd129;
	sample_rom[21][0] = 8'd130;
	sample_rom[21][1] = 8'd203;
	sample_rom[21][2] = 8'd243;
	sample_rom[21][3] = 8'd240;
	sample_rom[21][4] = 8'd196;
	sample_rom[21][5] = 8'd135;
	sample_rom[21][6] = 8'd82;
	sample_rom[21][7] = 8'd51;
	sample_rom[21][8] = 8'd54;
	sample_rom[21][9] = 8'd84;
	sample_rom[21][10] = 8'd130;
	sample_rom[21][11] = 8'd178;
	sample_rom[21][12] = 8'd213;
	sample_rom[21][13] = 8'd217;
	sample_rom[21][14] = 8'd196;
	sample_rom[21][15] = 8'd154;
	sample_rom[21][16] = 8'd116;
	sample_rom[21][17] = 8'd93;
	sample_rom[21][18] = 8'd94;
	sample_rom[21][19] = 8'd113;
	sample_rom[21][20] = 8'd140;
	sample_rom[21][21] = 8'd167;
	sample_rom[21][22] = 8'd187;
	sample_rom[21][23] = 8'd188;
	sample_rom[21][24] = 8'd177;
	sample_rom[21][25] = 8'd153;
	sample_rom[21][26] = 8'd130;
	sample_rom[21][27] = 8'd114;
	sample_rom[21][28] = 8'd117;
	sample_rom[21][29] = 8'd131;
	sample_rom[21][30] = 8'd150;
	sample_rom[21][31] = 8'd166;
	sample_rom[21][32] = 8'd174;
	sample_rom[21][33] = 8'd170;
	sample_rom[21][34] = 8'd156;
	sample_rom[21][35] = 8'd134;
	sample_rom[21][36] = 8'd121;
	sample_rom[21][37] = 8'd114;
	sample_rom[21][38] = 8'd117;
	sample_rom[21][39] = 8'd132;
	sample_rom[21][40] = 8'd150;
	sample_rom[21][41] = 8'd164;
	sample_rom[21][42] = 8'd169;
	sample_rom[21][43] = 8'd161;
	sample_rom[21][44] = 8'd145;
	sample_rom[21][45] = 8'd127;
	sample_rom[21][46] = 8'd113;
	sample_rom[21][47] = 8'd108;
	sample_rom[21][48] = 8'd112;
	sample_rom[21][49] = 8'd128;
	sample_rom[21][50] = 8'd146;
	sample_rom[21][51] = 8'd157;
	sample_rom[21][52] = 8'd160;
	sample_rom[21][53] = 8'd154;
	sample_rom[21][54] = 8'd137;
	sample_rom[21][55] = 8'd117;
	sample_rom[21][56] = 8'd109;
	sample_rom[21][57] = 8'd103;
	sample_rom[21][58] = 8'd114;
	sample_rom[21][59] = 8'd125;
	sample_rom[21][60] = 8'd139;
	sample_rom[21][61] = 8'd147;
	sample_rom[21][62] = 8'd148;
	sample_rom[21][63] = 8'd142;
	sample_rom[22][0] = 8'd129;
	sample_rom[22][1] = 8'd186;
	sample_rom[22][2] = 8'd221;
	sample_rom[22][3] = 8'd227;
	sample_rom[22][4] = 8'd209;
	sample_rom[22][5] = 8'd172;
	sample_rom[22][6] = 8'd134;
	sample_rom[22][7] = 8'd99;
	sample_rom[22][8] = 8'd82;
	sample_rom[22][9] = 8'd73;
	sample_rom[22][10] = 8'd88;
	sample_rom[22][11] = 8'd109;
	sample_rom[22][12] = 8'd142;
	sample_rom[22][13] = 8'd168;
	sample_rom[22][14] = 8'd184;
	sample_rom[22][15] = 8'd184;
	sample_rom[22][16] = 8'd170;
	sample_rom[22][17] = 8'd147;
	sample_rom[22][18] = 8'd121;
	sample_rom[22][19] = 8'd97;
	sample_rom[22][20] = 8'd88;
	sample_rom[22][21] = 8'd91;
	sample_rom[22][22] = 8'd103;
	sample_rom[22][23] = 8'd123;
	sample_rom[22][24] = 8'd149;
	sample_rom[22][25] = 8'd166;
	sample_rom[22][26] = 8'd170;
	sample_rom[22][27] = 8'd164;
	sample_rom[22][28] = 8'd151;
	sample_rom[22][29] = 8'd131;
	sample_rom[22][30] = 8'd112;
	sample_rom[22][31] = 8'd99;
	sample_rom[22][32] = 8'd97;
	sample_rom[22][33] = 8'd107;
	sample_rom[22][34] = 8'd120;
	sample_rom[22][35] = 8'd136;
	sample_rom[22][36] = 8'd149;
	sample_rom[22][37] = 8'd154;
	sample_rom[22][38] = 8'd152;
	sample_rom[22][39] = 8'd148;
	sample_rom[22][40] = 8'd137;
	sample_rom[22][41] = 8'd125;
	sample_rom[22][42] = 8'd122;
	sample_rom[22][43] = 8'd113;
	sample_rom[22][44] = 8'd115;
	sample_rom[22][45] = 8'd121;
	sample_rom[22][46] = 8'd125;
	sample_rom[22][47] = 8'd132;
	sample_rom[22][48] = 8'd136;
	sample_rom[22][49] = 8'd139;
	sample_rom[22][50] = 8'd139;
	sample_rom[22][51] = 8'd139;
	sample_rom[22][52] = 8'd137;
	sample_rom[22][53] = 8'd126;
	sample_rom[22][54] = 8'd118;
	sample_rom[22][55] = 8'd117;
	sample_rom[22][56] = 8'd118;
	sample_rom[22][57] = 8'd120;
	sample_rom[22][58] = 8'd127;
	sample_rom[22][59] = 8'd133;
	sample_rom[22][60] = 8'd138;
	sample_rom[22][61] = 8'd143;
	sample_rom[22][62] = 8'd141;
	sample_rom[22][63] = 8'd135;
	sample_rom[23][0] = 8'd130;
	sample_rom[23][1] = 8'd180;
	sample_rom[23][2] = 8'd218;
	sample_rom[23][3] = 8'd237;
	sample_rom[23][4] = 8'd237;
	sample_rom[23][5] = 8'd220;
	sample_rom[23][6] = 8'd190;
	sample_rom[23][7] = 8'd155;
	sample_rom[23][8] = 8'd118;
	sample_rom[23][9] = 8'd89;
	sample_rom[23][10] = 8'd67;
	sample_rom[23][11] = 8'd61;
	sample_rom[23][12] = 8'd70;
	sample_rom[23][13] = 8'd89;
	sample_rom[23][14] = 8'd117;
	sample_rom[23][15] = 8'd147;
	sample_rom[23][16] = 8'd173;
	sample_rom[23][17] = 8'd190;
	sample_rom[23][18] = 8'd195;
	sample_rom[23][19] = 8'd190;
	sample_rom[23][20] = 8'd173;
	sample_rom[23][21] = 8'd152;
	sample_rom[23][22] = 8'd129;
	sample_rom[23][23] = 8'd105;
	sample_rom[23][24] = 8'd92;
	sample_rom[23][25] = 8'd86;
	sample_rom[23][26] = 8'd90;
	sample_rom[23][27] = 8'd101;
	sample_rom[23][28] = 8'd120;
	sample_rom[23][29] = 8'd141;
	sample_rom[23][30] = 8'd155;
	sample_rom[23][31] = 8'd167;
	sample_rom[23][32] = 8'd173;
	sample_rom[23][33] = 8'd168;
	sample_rom[23][34] = 8'd155;
	sample_rom[23][35] = 8'd141;
	sample_rom[23][36] = 8'd123;
	sample_rom[23][37] = 8'd107;
	sample_rom[23][38] = 8'd101;
	sample_rom[23][39] = 8'd101;
	sample_rom[23][40] = 8'd106;
	sample_rom[23][41] = 8'd116;
	sample_rom[23][42] = 8'd127;
	sample_rom[23][43] = 8'd140;
	sample_rom[23][44] = 8'd151;
	sample_rom[23][45] = 8'd155;
	sample_rom[23][46] = 8'd157;
	sample_rom[23][47] = 8'd153;
	sample_rom[23][48] = 8'd144;
	sample_rom[23][49] = 8'd134;
	sample_rom[23][50] = 8'd123;
	sample_rom[23][51] = 8'd117;
	sample_rom[23][52] = 8'd112;
	sample_rom[23][53] = 8'd110;
	sample_rom[23][54] = 8'd111;
	sample_rom[23][55] = 8'd116;
	sample_rom[23][56] = 8'd122;
	sample_rom[23][57] = 8'd134;
	sample_rom[23][58] = 8'd144;
	sample_rom[23][59] = 8'd143;
	sample_rom[23][60] = 8'd145;
	sample_rom[23][61] = 8'd140;
	sample_rom[23][62] = 8'd135;
	sample_rom[23][63] = 8'd129;
	sample_rom[24][0] = 8'd131;
	sample_rom[24][1] = 8'd160;
	sample_rom[24][2] = 8'd181;
	sample_rom[24][3] = 8'd204;
	sample_rom[24][4] = 8'd221;
	sample_rom[24][5] = 8'd233;
	sample_rom[24][6] = 8'd241;
	sample_rom[24][7] = 8'd242;
	sample_rom[24][8] = 8'd240;
	sample_rom[24][9] = 8'd235;
	sample_rom[24][10] = 8'd225;
	sample_rom[24][11] = 8'd214;
	sample_rom[24][12] = 8'd203;
	sample_rom[24][13] = 8'd191;
	sample_rom[24][14] = 8'd182;
	sample_rom[24][15] = 8'd174;
	sample_rom[24][16] = 8'd167;
	sample_rom[24][17] = 8'd162;
	sample_rom[24][18] = 8'd161;
	sample_rom[24][19] = 8'd160;
	sample_rom[24][20] = 8'd162;
	sample_rom[24][21] = 8'd165;
	sample_rom[24][22] = 8'd167;
	sample_rom[24][23] = 8'd170;
	sample_rom[24][24] = 8'd173;
	sample_rom[24][25] = 8'd171;
	sample_rom[24][26] = 8'd169;
	sample_rom[24][27] = 8'd166;
	sample_rom[24][28] = 8'd160;
	sample_rom[24][29] = 8'd153;
	sample_rom[24][30] = 8'd146;
	sample_rom[24][31] = 8'd136;
	sample_rom[24][32] = 8'd128;
	sample_rom[24][33] = 8'd120;
	sample_rom[24][34] = 8'd112;
	sample_rom[24][35] = 8'd107;
	sample_rom[24][36] = 8'd107;
	sample_rom[24][37] = 8'd107;
	sample_rom[24][38] = 8'd113;
	sample_rom[24][39] = 8'd119;
	sample_rom[24][40] = 8'd131;
	sample_rom[24][41] = 8'd143;
	sample_rom[24][42] = 8'd157;
	sample_rom[24][43] = 8'd168;
	sample_rom[24][44] = 8'd179;
	sample_rom[24][45] = 8'd188;
	sample_rom[24][46] = 8'd195;
	sample_rom[24][47] = 8'd197;
	sample_rom[24][48] = 8'd197;
	sample_rom[24][49] = 8'd190;
	sample_rom[24][50] = 8'd183;
	sample_rom[24][51] = 8'd172;
	sample_rom[24][52] = 8'd160;
	sample_rom[24][53] = 8'd149;
	sample_rom[24][54] = 8'd136;
	sample_rom[24][55] = 8'd125;
	sample_rom[24][56] = 8'd113;
	sample_rom[24][57] = 8'd109;
	sample_rom[24][58] = 8'd105;
	sample_rom[24][59] = 8'd103;
	sample_rom[24][60] = 8'd105;
	sample_rom[24][61] = 8'd109;
	sample_rom[24][62] = 8'd113;
	sample_rom[24][63] = 8'd120;
	sample_rom[25][0] = 8'd131;
	sample_rom[25][1] = 8'd164;
	sample_rom[25][2] = 8'd191;
	sample_rom[25][3] = 8'd216;
	sample_rom[25][4] = 8'd233;
	sample_rom[25][5] = 8'd243;
	sample_rom[25][6] = 8'd246;
	sample_rom[25][7] = 8'd239;
	sample_rom[25][8] = 8'd231;
	sample_rom[25][9] = 8'd214;
	sample_rom[25][10] = 8'd194;
	sample_rom[25][11] = 8'd174;
	sample_rom[25][12] = 8'd154;
	sample_rom[25][13] = 8'd129;
	sample_rom[25][14] = 8'd110;
	sample_rom[25][15] = 8'd95;
	sample_rom[25][16] = 8'd83;
	sample_rom[25][17] = 8'd73;
	sample_rom[25][18] = 8'd73;
	sample_rom[25][19] = 8'd74;
	sample_rom[25][20] = 8'd83;
	sample_rom[25][21] = 8'd93;
	sample_rom[25][22] = 8'd107;
	sample_rom[25][23] = 8'd121;
	sample_rom[25][24] = 8'd138;
	sample_rom[25][25] = 8'd153;
	sample_rom[25][26] = 8'd163;
	sample_rom[25][27] = 8'd174;
	sample_rom[25][28] = 8'd184;
	sample_rom[25][29] = 8'd187;
	sample_rom[25][30] = 8'd188;
	sample_rom[25][31] = 8'd189;
	sample_rom[25][32] = 8'd185;
	sample_rom[25][33] = 8'd178;
	sample_rom[25][34] = 8'd169;
	sample_rom[25][35] = 8'd160;
	sample_rom[25][36] = 8'd152;
	sample_rom[25][37] = 8'd141;
	sample_rom[25][38] = 8'd134;
	sample_rom[25][39] = 8'd127;
	sample_rom[25][40] = 8'd122;
	sample_rom[25][41] = 8'd119;
	sample_rom[25][42] = 8'd117;
	sample_rom[25][43] = 8'd118;
	sample_rom[25][44] = 8'd119;
	sample_rom[25][45] = 8'd122;
	sample_rom[25][46] = 8'd125;
	sample_rom[25][47] = 8'd132;
	sample_rom[25][48] = 8'd137;
	sample_rom[25][49] = 8'd140;
	sample_rom[25][50] = 8'd144;
	sample_rom[25][51] = 8'd146;
	sample_rom[25][52] = 8'd147;
	sample_rom[25][53] = 8'd145;
	sample_rom[25][54] = 8'd144;
	sample_rom[25][55] = 8'd140;
	sample_rom[25][56] = 8'd139;
	sample_rom[25][57] = 8'd137;
	sample_rom[25][58] = 8'd135;
	sample_rom[25][59] = 8'd136;
	sample_rom[25][60] = 8'd134;
	sample_rom[25][61] = 8'd134;
	sample_rom[25][62] = 8'd132;
	sample_rom[25][63] = 8'd132;
	sample_rom[26][0] = 8'd130;
	sample_rom[26][1] = 8'd154;
	sample_rom[26][2] = 8'd175;
	sample_rom[26][3] = 8'd190;
	sample_rom[26][4] = 8'd206;
	sample_rom[26][5] = 8'd215;
	sample_rom[26][6] = 8'd219;
	sample_rom[26][7] = 8'd219;
	sample_rom[26][8] = 8'd218;
	sample_rom[26][9] = 8'd210;
	sample_rom[26][10] = 8'd201;
	sample_rom[26][11] = 8'd190;
	sample_rom[26][12] = 8'd177;
	sample_rom[26][13] = 8'd164;
	sample_rom[26][14] = 8'd152;
	sample_rom[26][15] = 8'd140;
	sample_rom[26][16] = 8'd126;
	sample_rom[26][17] = 8'd114;
	sample_rom[26][18] = 8'd104;
	sample_rom[26][19] = 8'd98;
	sample_rom[26][20] = 8'd95;
	sample_rom[26][21] = 8'd96;
	sample_rom[26][22] = 8'd98;
	sample_rom[26][23] = 8'd106;
	sample_rom[26][24] = 8'd112;
	sample_rom[26][25] = 8'd123;
	sample_rom[26][26] = 8'd131;
	sample_rom[26][27] = 8'd140;
	sample_rom[26][28] = 8'd147;
	sample_rom[26][29] = 8'd153;
	sample_rom[26][30] = 8'd157;
	sample_rom[26][31] = 8'd158;
	sample_rom[26][32] = 8'd160;
	sample_rom[26][33] = 8'd160;
	sample_rom[26][34] = 8'd160;
	sample_rom[26][35] = 8'd160;
	sample_rom[26][36] = 8'd160;
	sample_rom[26][37] = 8'd160;
	sample_rom[26][38] = 8'd159;
	sample_rom[26][39] = 8'd158;
	sample_rom[26][40] = 8'd155;
	sample_rom[26][41] = 8'd153;
	sample_rom[26][42] = 8'd150;
	sample_rom[26][43] = 8'd146;
	sample_rom[26][44] = 8'd145;
	sample_rom[26][45] = 8'd143;
	sample_rom[26][46] = 8'd141;
	sample_rom[26][47] = 8'd140;
	sample_rom[26][48] = 8'd136;
	sample_rom[26][49] = 8'd136;
	sample_rom[26][50] = 8'd135;
	sample_rom[26][51] = 8'd130;
	sample_rom[26][52] = 8'd126;
	sample_rom[26][53] = 8'd123;
	sample_rom[26][54] = 8'd121;
	sample_rom[26][55] = 8'd115;
	sample_rom[26][56] = 8'd113;
	sample_rom[26][57] = 8'd112;
	sample_rom[26][58] = 8'd113;
	sample_rom[26][59] = 8'd113;
	sample_rom[26][60] = 8'd113;
	sample_rom[26][61] = 8'd117;
	sample_rom[26][62] = 8'd121;
	sample_rom[26][63] = 8'd123;
	sample_rom[27][0] = 8'd131;
	sample_rom[27][1] = 8'd146;
	sample_rom[27][2] = 8'd159;
	sample_rom[27][3] = 8'd171;
	sample_rom[27][4] = 8'd181;
	sample_rom[27][5] = 8'd194;
	sample_rom[27][6] = 8'd204;
	sample_rom[27][7] = 8'd212;
	sample_rom[27][8] = 8'd220;
	sample_rom[27][9] = 8'd226;
	sample_rom[27][10] = 8'd232;
	sample_rom[27][11] = 8'd235;
	sample_rom[27][12] = 8'd238;
	sample_rom[27][13] = 8'd238;
	sample_rom[27][14] = 8'd238;
	sample_rom[27][15] = 8'd238;
	sample_rom[27][16] = 8'd235;
	sample_rom[27][17] = 8'd230;
	sample_rom[27][18] = 8'd226;
	sample_rom[27][19] = 8'd222;
	sample_rom[27][20] = 8'd217;
	sample_rom[27][21] = 8'd212;
	sample_rom[27][22] = 8'd205;
	sample_rom[27][23] = 8'd200;
	sample_rom[27][24] = 8'd194;
	sample_rom[27][25] = 8'd188;
	sample_rom[27][26] = 8'd183;
	sample_rom[27][27] = 8'd178;
	sample_rom[27][28] = 8'd172;
	sample_rom[27][29] = 8'd167;
	sample_rom[27][30] = 8'd165;
	sample_rom[27][31] = 8'd160;
	sample_rom[27][32] = 8'd158;
	sample_rom[27][33] = 8'd155;
	sample_rom[27][34] = 8'd152;
	sample_rom[27][35] = 8'd151;
	sample_rom[27][36] = 8'd149;
	sample_rom[27][37] = 8'd146;
	sample_rom[27][38] = 8'd145;
	sample_rom[27][39] = 8'd143;
	sample_rom[27][40] = 8'd142;
	sample_rom[27][41] = 8'd140;
	sample_rom[27][42] = 8'd139;
	sample_rom[27][43] = 8'd136;
	sample_rom[27][44] = 8'd135;
	sample_rom[27][45] = 8'd132;
	sample_rom[27][46] = 8'd131;
	sample_rom[27][47] = 8'd129;
	sample_rom[27][48] = 8'd129;
	sample_rom[27][49] = 8'd126;
	sample_rom[27][50] = 8'd124;
	sample_rom[27][51] = 8'd123;
	sample_rom[27][52] = 8'd123;
	sample_rom[27][53] = 8'd121;
	sample_rom[27][54] = 8'd120;
	sample_rom[27][55] = 8'd119;
	sample_rom[27][56] = 8'd118;
	sample_rom[27][57] = 8'd120;
	sample_rom[27][58] = 8'd121;
	sample_rom[27][59] = 8'd122;
	sample_rom[27][60] = 8'd123;
	sample_rom[27][61] = 8'd124;
	sample_rom[27][62] = 8'd124;
	sample_rom[27][63] = 8'd126;
	sample_rom[28][0] = 8'd130;
	sample_rom[28][1] = 8'd141;
	sample_rom[28][2] = 8'd151;
	sample_rom[28][3] = 8'd158;
	sample_rom[28][4] = 8'd167;
	sample_rom[28][5] = 8'd175;
	sample_rom[28][6] = 8'd182;
	sample_rom[28][7] = 8'd191;
	sample_rom[28][8] = 8'd195;
	sample_rom[28][9] = 8'd201;
	sample_rom[28][10] = 8'd203;
	sample_rom[28][11] = 8'd207;
	sample_rom[28][12] = 8'd210;
	sample_rom[28][13] = 8'd211;
	sample_rom[28][14] = 8'd210;
	sample_rom[28][15] = 8'd211;
	sample_rom[28][16] = 8'd208;
	sample_rom[28][17] = 8'd205;
	sample_rom[28][18] = 8'd203;
	sample_rom[28][19] = 8'd198;
	sample_rom[28][20] = 8'd193;
	sample_rom[28][21] = 8'd189;
	sample_rom[28][22] = 8'd183;
	sample_rom[28][23] = 8'd177;
	sample_rom[28][24] = 8'd172;
	sample_rom[28][25] = 8'd164;
	sample_rom[28][26] = 8'd159;
	sample_rom[28][27] = 8'd153;
	sample_rom[28][28] = 8'd145;
	sample_rom[28][29] = 8'd139;
	sample_rom[28][30] = 8'd135;
	sample_rom[28][31] = 8'd129;
	sample_rom[28][32] = 8'd123;
	sample_rom[28][33] = 8'd118;
	sample_rom[28][34] = 8'd113;
	sample_rom[28][35] = 8'd109;
	sample_rom[28][36] = 8'd106;
	sample_rom[28][37] = 8'd100;
	sample_rom[28][38] = 8'd98;
	sample_rom[28][39] = 8'd96;
	sample_rom[28][40] = 8'd94;
	sample_rom[28][41] = 8'd92;
	sample_rom[28][42] = 8'd91;
	sample_rom[28][43] = 8'd89;
	sample_rom[28][44] = 8'd89;
	sample_rom[28][45] = 8'd88;
	sample_rom[28][46] = 8'd88;
	sample_rom[28][47] = 8'd88;
	sample_rom[28][48] = 8'd89;
	sample_rom[28][49] = 8'd89;
	sample_rom[28][50] = 8'd90;
	sample_rom[28][51] = 8'd91;
	sample_rom[28][52] = 8'd93;
	sample_rom[28][53] = 8'd94;
	sample_rom[28][54] = 8'd97;
	sample_rom[28][55] = 8'd99;
	sample_rom[28][56] = 8'd101;
	sample_rom[28][57] = 8'd104;
	sample_rom[28][58] = 8'd107;
	sample_rom[28][59] = 8'd111;
	sample_rom[28][60] = 8'd114;
	sample_rom[28][61] = 8'd119;
	sample_rom[28][62] = 8'd121;
	sample_rom[28][63] = 8'd124;
	sample_rom[29][0] = 8'd131;
	sample_rom[29][1] = 8'd140;
	sample_rom[29][2] = 8'd151;
	sample_rom[29][3] = 8'd159;
	sample_rom[29][4] = 8'd166;
	sample_rom[29][5] = 8'd174;
	sample_rom[29][6] = 8'd183;
	sample_rom[29][7] = 8'd190;
	sample_rom[29][8] = 8'd197;
	sample_rom[29][9] = 8'd204;
	sample_rom[29][10] = 8'd210;
	sample_rom[29][11] = 8'd216;
	sample_rom[29][12] = 8'd221;
	sample_rom[29][13] = 8'd225;
	sample_rom[29][14] = 8'd230;
	sample_rom[29][15] = 8'd233;
	sample_rom[29][16] = 8'd235;
	sample_rom[29][17] = 8'd238;
	sample_rom[29][18] = 8'd239;
	sample_rom[29][19] = 8'd241;
	sample_rom[29][20] = 8'd240;
	sample_rom[29][21] = 8'd241;
	sample_rom[29][22] = 8'd239;
	sample_rom[29][23] = 8'd240;
	sample_rom[29][24] = 8'd238;
	sample_rom[29][25] = 8'd236;
	sample_rom[29][26] = 8'd233;
	sample_rom[29][27] = 8'd230;
	sample_rom[29][28] = 8'd228;
	sample_rom[29][29] = 8'd225;
	sample_rom[29][30] = 8'd223;
	sample_rom[29][31] = 8'd219;
	sample_rom[29][32] = 8'd215;
	sample_rom[29][33] = 8'd211;
	sample_rom[29][34] = 8'd206;
	sample_rom[29][35] = 8'd203;
	sample_rom[29][36] = 8'd199;
	sample_rom[29][37] = 8'd195;
	sample_rom[29][38] = 8'd191;
	sample_rom[29][39] = 8'd187;
	sample_rom[29][40] = 8'd183;
	sample_rom[29][41] = 8'd179;
	sample_rom[29][42] = 8'd177;
	sample_rom[29][43] = 8'd171;
	sample_rom[29][44] = 8'd170;
	sample_rom[29][45] = 8'd167;
	sample_rom[29][46] = 8'd163;
	sample_rom[29][47] = 8'd160;
	sample_rom[29][48] = 8'd158;
	sample_rom[29][49] = 8'd156;
	sample_rom[29][50] = 8'd153;
	sample_rom[29][51] = 8'd151;
	sample_rom[29][52] = 8'd148;
	sample_rom[29][53] = 8'd146;
	sample_rom[29][54] = 8'd144;
	sample_rom[29][55] = 8'd143;
	sample_rom[29][56] = 8'd139;
	sample_rom[29][57] = 8'd138;
	sample_rom[29][58] = 8'd137;
	sample_rom[29][59] = 8'd135;
	sample_rom[29][60] = 8'd134;
	sample_rom[29][61] = 8'd132;
	sample_rom[29][62] = 8'd128;
	sample_rom[29][63] = 8'd128;
	sample_rom[30][0] = 8'd132;
	sample_rom[30][1] = 8'd140;
	sample_rom[30][2] = 8'd149;
	sample_rom[30][3] = 8'd156;
	sample_rom[30][4] = 8'd164;
	sample_rom[30][5] = 8'd170;
	sample_rom[30][6] = 8'd178;
	sample_rom[30][7] = 8'd186;
	sample_rom[30][8] = 8'd192;
	sample_rom[30][9] = 8'd199;
	sample_rom[30][10] = 8'd206;
	sample_rom[30][11] = 8'd212;
	sample_rom[30][12] = 8'd217;
	sample_rom[30][13] = 8'd223;
	sample_rom[30][14] = 8'd227;
	sample_rom[30][15] = 8'd232;
	sample_rom[30][16] = 8'd236;
	sample_rom[30][17] = 8'd240;
	sample_rom[30][18] = 8'd241;
	sample_rom[30][19] = 8'd244;
	sample_rom[30][20] = 8'd246;
	sample_rom[30][21] = 8'd248;
	sample_rom[30][22] = 8'd248;
	sample_rom[30][23] = 8'd250;
	sample_rom[30][24] = 8'd250;
	sample_rom[30][25] = 8'd251;
	sample_rom[30][26] = 8'd249;
	sample_rom[30][27] = 8'd249;
	sample_rom[30][28] = 8'd248;
	sample_rom[30][29] = 8'd245;
	sample_rom[30][30] = 8'd244;
	sample_rom[30][31] = 8'd241;
	sample_rom[30][32] = 8'd238;
	sample_rom[30][33] = 8'd236;
	sample_rom[30][34] = 8'd232;
	sample_rom[30][35] = 8'd230;
	sample_rom[30][36] = 8'd226;
	sample_rom[30][37] = 8'd223;
	sample_rom[30][38] = 8'd219;
	sample_rom[30][39] = 8'd214;
	sample_rom[30][40] = 8'd210;
	sample_rom[30][41] = 8'd206;
	sample_rom[30][42] = 8'd203;
	sample_rom[30][43] = 8'd198;
	sample_rom[30][44] = 8'd194;
	sample_rom[30][45] = 8'd190;
	sample_rom[30][46] = 8'd188;
	sample_rom[30][47] = 8'd183;
	sample_rom[30][48] = 8'd179;
	sample_rom[30][49] = 8'd175;
	sample_rom[30][50] = 8'd171;
	sample_rom[30][51] = 8'd166;
	sample_rom[30][52] = 8'd164;
	sample_rom[30][53] = 8'd160;
	sample_rom[30][54] = 8'd157;
	sample_rom[30][55] = 8'd153;
	sample_rom[30][56] = 8'd150;
	sample_rom[30][57] = 8'd146;
	sample_rom[30][58] = 8'd144;
	sample_rom[30][59] = 8'd142;
	sample_rom[30][60] = 8'd138;
	sample_rom[30][61] = 8'd136;
	sample_rom[30][62] = 8'd131;
	sample_rom[30][63] = 8'd129;
	sample_rom[31][0] = 8'd128;
	sample_rom[31][1] = 8'd128;
	sample_rom[31][2] = 8'd128;
	sample_rom[31][3] = 8'd128;
	sample_rom[31][4] = 8'd128;
	sample_rom[31][5] = 8'd128;
	sample_rom[31][6] = 8'd128;
	sample_rom[31][7] = 8'd128;
	sample_rom[31][8] = 8'd128;
	sample_rom[31][9] = 8'd128;
	sample_rom[31][10] = 8'd128;
	sample_rom[31][11] = 8'd128;
	sample_rom[31][12] = 8'd128;
	sample_rom[31][13] = 8'd128;
	sample_rom[31][14] = 8'd128;
	sample_rom[31][15] = 8'd128;
	sample_rom[31][16] = 8'd128;
	sample_rom[31][17] = 8'd128;
	sample_rom[31][18] = 8'd128;
	sample_rom[31][19] = 8'd128;
	sample_rom[31][20] = 8'd128;
	sample_rom[31][21] = 8'd128;
	sample_rom[31][22] = 8'd128;
	sample_rom[31][23] = 8'd128;
	sample_rom[31][24] = 8'd128;
	sample_rom[31][25] = 8'd128;
	sample_rom[31][26] = 8'd128;
	sample_rom[31][27] = 8'd128;
	sample_rom[31][28] = 8'd128;
	sample_rom[31][29] = 8'd128;
	sample_rom[31][30] = 8'd128;
	sample_rom[31][31] = 8'd128;
	sample_rom[31][32] = 8'd128;
	sample_rom[31][33] = 8'd128;
	sample_rom[31][34] = 8'd128;
	sample_rom[31][35] = 8'd128;
	sample_rom[31][36] = 8'd128;
	sample_rom[31][37] = 8'd128;
	sample_rom[31][38] = 8'd128;
	sample_rom[31][39] = 8'd128;
	sample_rom[31][40] = 8'd128;
	sample_rom[31][41] = 8'd128;
	sample_rom[31][42] = 8'd128;
	sample_rom[31][43] = 8'd128;
	sample_rom[31][44] = 8'd128;
	sample_rom[31][45] = 8'd128;
	sample_rom[31][46] = 8'd128;
	sample_rom[31][47] = 8'd128;
	sample_rom[31][48] = 8'd128;
	sample_rom[31][49] = 8'd128;
	sample_rom[31][50] = 8'd128;
	sample_rom[31][51] = 8'd128;
	sample_rom[31][52] = 8'd128;
	sample_rom[31][53] = 8'd128;
	sample_rom[31][54] = 8'd128;
	sample_rom[31][55] = 8'd128;
	sample_rom[31][56] = 8'd128;
	sample_rom[31][57] = 8'd128;
	sample_rom[31][58] = 8'd128;
	sample_rom[31][59] = 8'd128;
	sample_rom[31][60] = 8'd128;
	sample_rom[31][61] = 8'd128;
	sample_rom[31][62] = 8'd128;
	sample_rom[31][63] = 8'd128;
	sample_rom[32][0] = 8'd131;
	sample_rom[32][1] = 8'd137;
	sample_rom[32][2] = 8'd144;
	sample_rom[32][3] = 8'd150;
	sample_rom[32][4] = 8'd156;
	sample_rom[32][5] = 8'd160;
	sample_rom[32][6] = 8'd164;
	sample_rom[32][7] = 8'd170;
	sample_rom[32][8] = 8'd175;
	sample_rom[32][9] = 8'd181;
	sample_rom[32][10] = 8'd187;
	sample_rom[32][11] = 8'd192;
	sample_rom[32][12] = 8'd197;
	sample_rom[32][13] = 8'd202;
	sample_rom[32][14] = 8'd207;
	sample_rom[32][15] = 8'd212;
	sample_rom[32][16] = 8'd216;
	sample_rom[32][17] = 8'd220;
	sample_rom[32][18] = 8'd222;
	sample_rom[32][19] = 8'd224;
	sample_rom[32][20] = 8'd227;
	sample_rom[32][21] = 8'd231;
	sample_rom[32][22] = 8'd233;
	sample_rom[32][23] = 8'd236;
	sample_rom[32][24] = 8'd238;
	sample_rom[32][25] = 8'd241;
	sample_rom[32][26] = 8'd242;
	sample_rom[32][27] = 8'd244;
	sample_rom[32][28] = 8'd245;
	sample_rom[32][29] = 8'd246;
	sample_rom[32][30] = 8'd247;
	sample_rom[32][31] = 8'd247;
	sample_rom[32][32] = 8'd247;
	sample_rom[32][33] = 8'd247;
	sample_rom[32][34] = 8'd246;
	sample_rom[32][35] = 8'd245;
	sample_rom[32][36] = 8'd244;
	sample_rom[32][37] = 8'd242;
	sample_rom[32][38] = 8'd241;
	sample_rom[32][39] = 8'd238;
	sample_rom[32][40] = 8'd236;
	sample_rom[32][41] = 8'd233;
	sample_rom[32][42] = 8'd231;
	sample_rom[32][43] = 8'd227;
	sample_rom[32][44] = 8'd224;
	sample_rom[32][45] = 8'd222;
	sample_rom[32][46] = 8'd220;
	sample_rom[32][47] = 8'd216;
	sample_rom[32][48] = 8'd212;
	sample_rom[32][49] = 8'd207;
	sample_rom[32][50] = 8'd202;
	sample_rom[32][51] = 8'd197;
	sample_rom[32][52] = 8'd192;
	sample_rom[32][53] = 8'd187;
	sample_rom[32][54] = 8'd181;
	sample_rom[32][55] = 8'd175;
	sample_rom[32][56] = 8'd170;
	sample_rom[32][57] = 8'd164;
	sample_rom[32][58] = 8'd160;
	sample_rom[32][59] = 8'd156;
	sample_rom[32][60] = 8'd150;
	sample_rom[32][61] = 8'd144;
	sample_rom[32][62] = 8'd137;
	sample_rom[32][63] = 8'd131;
	sample_rom[33][0] = 8'd131;
	sample_rom[33][1] = 8'd152;
	sample_rom[33][2] = 8'd172;
	sample_rom[33][3] = 8'd188;
	sample_rom[33][4] = 8'd199;
	sample_rom[33][5] = 8'd206;
	sample_rom[33][6] = 8'd206;
	sample_rom[33][7] = 8'd200;
	sample_rom[33][8] = 8'd190;
	sample_rom[33][9] = 8'd174;
	sample_rom[33][10] = 8'd158;
	sample_rom[33][11] = 8'd139;
	sample_rom[33][12] = 8'd121;
	sample_rom[33][13] = 8'd105;
	sample_rom[33][14] = 8'd95;
	sample_rom[33][15] = 8'd89;
	sample_rom[33][16] = 8'd87;
	sample_rom[33][17] = 8'd91;
	sample_rom[33][18] = 8'd101;
	sample_rom[33][19] = 8'd115;
	sample_rom[33][20] = 8'd134;
	sample_rom[33][21] = 8'd155;
	sample_rom[33][22] = 8'd175;
	sample_rom[33][23] = 8'd194;
	sample_rom[33][24] = 8'd212;
	sample_rom[33][25] = 8'd223;
	sample_rom[33][26] = 8'd229;
	sample_rom[33][27] = 8'd231;
	sample_rom[33][28] = 8'd225;
	sample_rom[33][29] = 8'd216;
	sample_rom[33][30] = 8'd201;
	sample_rom[33][31] = 8'd182;
	sample_rom[33][32] = 8'd162;
	sample_rom[33][33] = 8'd144;
	sample_rom[33][34] = 8'd124;
	sample_rom[33][35] = 8'd110;
	sample_rom[33][36] = 8'd100;
	sample_rom[33][37] = 8'd95;
	sample_rom[33][38] = 8'd97;
	sample_rom[33][39] = 8'd102;
	sample_rom[33][40] = 8'd113;
	sample_rom[33][41] = 8'd129;
	sample_rom[33][42] = 8'd148;
	sample_rom[33][43] = 8'd167;
	sample_rom[33][44] = 8'd185;
	sample_rom[33][45] = 8'd202;
	sample_rom[33][46] = 8'd213;
	sample_rom[33][47] = 8'd220;
	sample_rom[33][48] = 8'd222;
	sample_rom[33][49] = 8'd217;
	sample_rom[33][50] = 8'd206;
	sample_rom[33][51] = 8'd191;
	sample_rom[33][52] = 8'd172;
	sample_rom[33][53] = 8'd151;
	sample_rom[33][54] = 8'd128;
	sample_rom[33][55] = 8'd109;
	sample_rom[33][56] = 8'd91;
	sample_rom[33][57] = 8'd79;
	sample_rom[33][58] = 8'd71;
	sample_rom[33][59] = 8'd68;
	sample_rom[33][60] = 8'd73;
	sample_rom[33][61] = 8'd82;
	sample_rom[33][62] = 8'd95;
	sample_rom[33][63] = 8'd111;
	sample_rom[34][0] = 8'd131;
	sample_rom[34][1] = 8'd160;
	sample_rom[34][2] = 8'd181;
	sample_rom[34][3] = 8'd204;
	sample_rom[34][4] = 8'd221;
	sample_rom[34][5] = 8'd233;
	sample_rom[34][6] = 8'd241;
	sample_rom[34][7] = 8'd242;
	sample_rom[34][8] = 8'd240;
	sample_rom[34][9] = 8'd235;
	sample_rom[34][10] = 8'd225;
	sample_rom[34][11] = 8'd214;
	sample_rom[34][12] = 8'd203;
	sample_rom[34][13] = 8'd191;
	sample_rom[34][14] = 8'd182;
	sample_rom[34][15] = 8'd174;
	sample_rom[34][16] = 8'd167;
	sample_rom[34][17] = 8'd162;
	sample_rom[34][18] = 8'd161;
	sample_rom[34][19] = 8'd160;
	sample_rom[34][20] = 8'd162;
	sample_rom[34][21] = 8'd165;
	sample_rom[34][22] = 8'd167;
	sample_rom[34][23] = 8'd170;
	sample_rom[34][24] = 8'd173;
	sample_rom[34][25] = 8'd171;
	sample_rom[34][26] = 8'd169;
	sample_rom[34][27] = 8'd166;
	sample_rom[34][28] = 8'd160;
	sample_rom[34][29] = 8'd153;
	sample_rom[34][30] = 8'd146;
	sample_rom[34][31] = 8'd136;
	sample_rom[34][32] = 8'd128;
	sample_rom[34][33] = 8'd120;
	sample_rom[34][34] = 8'd112;
	sample_rom[34][35] = 8'd107;
	sample_rom[34][36] = 8'd107;
	sample_rom[34][37] = 8'd107;
	sample_rom[34][38] = 8'd113;
	sample_rom[34][39] = 8'd119;
	sample_rom[34][40] = 8'd131;
	sample_rom[34][41] = 8'd143;
	sample_rom[34][42] = 8'd157;
	sample_rom[34][43] = 8'd168;
	sample_rom[34][44] = 8'd179;
	sample_rom[34][45] = 8'd188;
	sample_rom[34][46] = 8'd195;
	sample_rom[34][47] = 8'd197;
	sample_rom[34][48] = 8'd197;
	sample_rom[34][49] = 8'd190;
	sample_rom[34][50] = 8'd183;
	sample_rom[34][51] = 8'd172;
	sample_rom[34][52] = 8'd160;
	sample_rom[34][53] = 8'd149;
	sample_rom[34][54] = 8'd136;
	sample_rom[34][55] = 8'd125;
	sample_rom[34][56] = 8'd113;
	sample_rom[34][57] = 8'd109;
	sample_rom[34][58] = 8'd105;
	sample_rom[34][59] = 8'd103;
	sample_rom[34][60] = 8'd105;
	sample_rom[34][61] = 8'd109;
	sample_rom[34][62] = 8'd113;
	sample_rom[34][63] = 8'd120;
	sample_rom[35][0] = 8'd128;
	sample_rom[35][1] = 8'd200;
	sample_rom[35][2] = 8'd238;
	sample_rom[35][3] = 8'd243;
	sample_rom[35][4] = 8'd222;
	sample_rom[35][5] = 8'd193;
	sample_rom[35][6] = 8'd172;
	sample_rom[35][7] = 8'd164;
	sample_rom[35][8] = 8'd164;
	sample_rom[35][9] = 8'd173;
	sample_rom[35][10] = 8'd180;
	sample_rom[35][11] = 8'd185;
	sample_rom[35][12] = 8'd180;
	sample_rom[35][13] = 8'd180;
	sample_rom[35][14] = 8'd189;
	sample_rom[35][15] = 8'd194;
	sample_rom[35][16] = 8'd205;
	sample_rom[35][17] = 8'd202;
	sample_rom[35][18] = 8'd195;
	sample_rom[35][19] = 8'd175;
	sample_rom[35][20] = 8'd157;
	sample_rom[35][21] = 8'd138;
	sample_rom[35][22] = 8'd132;
	sample_rom[35][23] = 8'd140;
	sample_rom[35][24] = 8'd151;
	sample_rom[35][25] = 8'd155;
	sample_rom[35][26] = 8'd145;
	sample_rom[35][27] = 8'd121;
	sample_rom[35][28] = 8'd101;
	sample_rom[35][29] = 8'd92;
	sample_rom[35][30] = 8'd93;
	sample_rom[35][31] = 8'd105;
	sample_rom[35][32] = 8'd127;
	sample_rom[35][33] = 8'd155;
	sample_rom[35][34] = 8'd166;
	sample_rom[35][35] = 8'd161;
	sample_rom[35][36] = 8'd147;
	sample_rom[35][37] = 8'd132;
	sample_rom[35][38] = 8'd127;
	sample_rom[35][39] = 8'd135;
	sample_rom[35][40] = 8'd149;
	sample_rom[35][41] = 8'd161;
	sample_rom[35][42] = 8'd164;
	sample_rom[35][43] = 8'd161;
	sample_rom[35][44] = 8'd148;
	sample_rom[35][45] = 8'd131;
	sample_rom[35][46] = 8'd118;
	sample_rom[35][47] = 8'd115;
	sample_rom[35][48] = 8'd119;
	sample_rom[35][49] = 8'd125;
	sample_rom[35][50] = 8'd133;
	sample_rom[35][51] = 8'd135;
	sample_rom[35][52] = 8'd140;
	sample_rom[35][53] = 8'd147;
	sample_rom[35][54] = 8'd154;
	sample_rom[35][55] = 8'd162;
	sample_rom[35][56] = 8'd160;
	sample_rom[35][57] = 8'd148;
	sample_rom[35][58] = 8'd121;
	sample_rom[35][59] = 8'd90;
	sample_rom[35][60] = 8'd67;
	sample_rom[35][61] = 8'd63;
	sample_rom[35][62] = 8'd76;
	sample_rom[35][63] = 8'd101;
	sample_rom[36][0] = 8'd128;
	sample_rom[36][1] = 8'd196;
	sample_rom[36][2] = 8'd232;
	sample_rom[36][3] = 8'd229;
	sample_rom[36][4] = 8'd202;
	sample_rom[36][5] = 8'd170;
	sample_rom[36][6] = 8'd146;
	sample_rom[36][7] = 8'd136;
	sample_rom[36][8] = 8'd139;
	sample_rom[36][9] = 8'd151;
	sample_rom[36][10] = 8'd162;
	sample_rom[36][11] = 8'd164;
	sample_rom[36][12] = 8'd156;
	sample_rom[36][13] = 8'd146;
	sample_rom[36][14] = 8'd142;
	sample_rom[36][15] = 8'd143;
	sample_rom[36][16] = 8'd151;
	sample_rom[36][17] = 8'd160;
	sample_rom[36][18] = 8'd165;
	sample_rom[36][19] = 8'd161;
	sample_rom[36][20] = 8'd150;
	sample_rom[36][21] = 8'd139;
	sample_rom[36][22] = 8'd131;
	sample_rom[36][23] = 8'd135;
	sample_rom[36][24] = 8'd139;
	sample_rom[36][25] = 8'd142;
	sample_rom[36][26] = 8'd139;
	sample_rom[36][27] = 8'd136;
	sample_rom[36][28] = 8'd126;
	sample_rom[36][29] = 8'd120;
	sample_rom[36][30] = 8'd120;
	sample_rom[36][31] = 8'd124;
	sample_rom[36][32] = 8'd133;
	sample_rom[36][33] = 8'd139;
	sample_rom[36][34] = 8'd134;
	sample_rom[36][35] = 8'd133;
	sample_rom[36][36] = 8'd128;
	sample_rom[36][37] = 8'd123;
	sample_rom[36][38] = 8'd125;
	sample_rom[36][39] = 8'd135;
	sample_rom[36][40] = 8'd143;
	sample_rom[36][41] = 8'd146;
	sample_rom[36][42] = 8'd140;
	sample_rom[36][43] = 8'd132;
	sample_rom[36][44] = 8'd125;
	sample_rom[36][45] = 8'd125;
	sample_rom[36][46] = 8'd131;
	sample_rom[36][47] = 8'd139;
	sample_rom[36][48] = 8'd146;
	sample_rom[36][49] = 8'd147;
	sample_rom[36][50] = 8'd141;
	sample_rom[36][51] = 8'd130;
	sample_rom[36][52] = 8'd127;
	sample_rom[36][53] = 8'd131;
	sample_rom[36][54] = 8'd142;
	sample_rom[36][55] = 8'd153;
	sample_rom[36][56] = 8'd161;
	sample_rom[36][57] = 8'd154;
	sample_rom[36][58] = 8'd131;
	sample_rom[36][59] = 8'd97;
	sample_rom[36][60] = 8'd67;
	sample_rom[36][61] = 8'd58;
	sample_rom[36][62] = 8'd71;
	sample_rom[36][63] = 8'd99;
	sample_rom[37][0] = 8'd131;
	sample_rom[37][1] = 8'd155;
	sample_rom[37][2] = 8'd177;
	sample_rom[37][3] = 8'd195;
	sample_rom[37][4] = 8'd212;
	sample_rom[37][5] = 8'd227;
	sample_rom[37][6] = 8'd239;
	sample_rom[37][7] = 8'd245;
	sample_rom[37][8] = 8'd250;
	sample_rom[37][9] = 8'd250;
	sample_rom[37][10] = 8'd247;
	sample_rom[37][11] = 8'd241;
	sample_rom[37][12] = 8'd235;
	sample_rom[37][13] = 8'd224;
	sample_rom[37][14] = 8'd216;
	sample_rom[37][15] = 8'd206;
	sample_rom[37][16] = 8'd196;
	sample_rom[37][17] = 8'd186;
	sample_rom[37][18] = 8'd177;
	sample_rom[37][19] = 8'd169;
	sample_rom[37][20] = 8'd162;
	sample_rom[37][21] = 8'd157;
	sample_rom[37][22] = 8'd151;
	sample_rom[37][23] = 8'd149;
	sample_rom[37][24] = 8'd145;
	sample_rom[37][25] = 8'd141;
	sample_rom[37][26] = 8'd138;
	sample_rom[37][27] = 8'd135;
	sample_rom[37][28] = 8'd131;
	sample_rom[37][29] = 8'd127;
	sample_rom[37][30] = 8'd122;
	sample_rom[37][31] = 8'd117;
	sample_rom[37][32] = 8'd115;
	sample_rom[37][33] = 8'd110;
	sample_rom[37][34] = 8'd105;
	sample_rom[37][35] = 8'd104;
	sample_rom[37][36] = 8'd102;
	sample_rom[37][37] = 8'd100;
	sample_rom[37][38] = 8'd100;
	sample_rom[37][39] = 8'd101;
	sample_rom[37][40] = 8'd103;
	sample_rom[37][41] = 8'd107;
	sample_rom[37][42] = 8'd111;
	sample_rom[37][43] = 8'd115;
	sample_rom[37][44] = 8'd120;
	sample_rom[37][45] = 8'd123;
	sample_rom[37][46] = 8'd128;
	sample_rom[37][47] = 8'd130;
	sample_rom[37][48] = 8'd131;
	sample_rom[37][49] = 8'd133;
	sample_rom[37][50] = 8'd134;
	sample_rom[37][51] = 8'd133;
	sample_rom[37][52] = 8'd132;
	sample_rom[37][53] = 8'd130;
	sample_rom[37][54] = 8'd129;
	sample_rom[37][55] = 8'd124;
	sample_rom[37][56] = 8'd123;
	sample_rom[37][57] = 8'd121;
	sample_rom[37][58] = 8'd121;
	sample_rom[37][59] = 8'd121;
	sample_rom[37][60] = 8'd121;
	sample_rom[37][61] = 8'd124;
	sample_rom[37][62] = 8'd123;
	sample_rom[37][63] = 8'd127;
	sample_rom[38][0] = 8'd131;
	sample_rom[38][1] = 8'd176;
	sample_rom[38][2] = 8'd213;
	sample_rom[38][3] = 8'd238;
	sample_rom[38][4] = 8'd248;
	sample_rom[38][5] = 8'd247;
	sample_rom[38][6] = 8'd234;
	sample_rom[38][7] = 8'd218;
	sample_rom[38][8] = 8'd200;
	sample_rom[38][9] = 8'd186;
	sample_rom[38][10] = 8'd180;
	sample_rom[38][11] = 8'd180;
	sample_rom[38][12] = 8'd186;
	sample_rom[38][13] = 8'd192;
	sample_rom[38][14] = 8'd193;
	sample_rom[38][15] = 8'd193;
	sample_rom[38][16] = 8'd182;
	sample_rom[38][17] = 8'd167;
	sample_rom[38][18] = 8'd148;
	sample_rom[38][19] = 8'd127;
	sample_rom[38][20] = 8'd110;
	sample_rom[38][21] = 8'd96;
	sample_rom[38][22] = 8'd91;
	sample_rom[38][23] = 8'd85;
	sample_rom[38][24] = 8'd89;
	sample_rom[38][25] = 8'd93;
	sample_rom[38][26] = 8'd96;
	sample_rom[38][27] = 8'd97;
	sample_rom[38][28] = 8'd97;
	sample_rom[38][29] = 8'd97;
	sample_rom[38][30] = 8'd99;
	sample_rom[38][31] = 8'd98;
	sample_rom[38][32] = 8'd105;
	sample_rom[38][33] = 8'd111;
	sample_rom[38][34] = 8'd120;
	sample_rom[38][35] = 8'd132;
	sample_rom[38][36] = 8'd139;
	sample_rom[38][37] = 8'd146;
	sample_rom[38][38] = 8'd149;
	sample_rom[38][39] = 8'd149;
	sample_rom[38][40] = 8'd145;
	sample_rom[38][41] = 8'd139;
	sample_rom[38][42] = 8'd133;
	sample_rom[38][43] = 8'd124;
	sample_rom[38][44] = 8'd118;
	sample_rom[38][45] = 8'd113;
	sample_rom[38][46] = 8'd108;
	sample_rom[38][47] = 8'd106;
	sample_rom[38][48] = 8'd106;
	sample_rom[38][49] = 8'd104;
	sample_rom[38][50] = 8'd105;
	sample_rom[38][51] = 8'd106;
	sample_rom[38][52] = 8'd109;
	sample_rom[38][53] = 8'd107;
	sample_rom[38][54] = 8'd110;
	sample_rom[38][55] = 8'd111;
	sample_rom[38][56] = 8'd112;
	sample_rom[38][57] = 8'd115;
	sample_rom[38][58] = 8'd114;
	sample_rom[38][59] = 8'd116;
	sample_rom[38][60] = 8'd117;
	sample_rom[38][61] = 8'd119;
	sample_rom[38][62] = 8'd121;
	sample_rom[38][63] = 8'd125;
	sample_rom[39][0] = 8'd132;
	sample_rom[39][1] = 8'd172;
	sample_rom[39][2] = 8'd206;
	sample_rom[39][3] = 8'd227;
	sample_rom[39][4] = 8'd232;
	sample_rom[39][5] = 8'd223;
	sample_rom[39][6] = 8'd203;
	sample_rom[39][7] = 8'd179;
	sample_rom[39][8] = 8'd157;
	sample_rom[39][9] = 8'd142;
	sample_rom[39][10] = 8'd137;
	sample_rom[39][11] = 8'd139;
	sample_rom[39][12] = 8'd152;
	sample_rom[39][13] = 8'd160;
	sample_rom[39][14] = 8'd167;
	sample_rom[39][15] = 8'd172;
	sample_rom[39][16] = 8'd169;
	sample_rom[39][17] = 8'd162;
	sample_rom[39][18] = 8'd154;
	sample_rom[39][19] = 8'd146;
	sample_rom[39][20] = 8'd147;
	sample_rom[39][21] = 8'd151;
	sample_rom[39][22] = 8'd160;
	sample_rom[39][23] = 8'd170;
	sample_rom[39][24] = 8'd180;
	sample_rom[39][25] = 8'd184;
	sample_rom[39][26] = 8'd184;
	sample_rom[39][27] = 8'd174;
	sample_rom[39][28] = 8'd159;
	sample_rom[39][29] = 8'd142;
	sample_rom[39][30] = 8'd127;
	sample_rom[39][31] = 8'd117;
	sample_rom[39][32] = 8'd116;
	sample_rom[39][33] = 8'd122;
	sample_rom[39][34] = 8'd132;
	sample_rom[39][35] = 8'd144;
	sample_rom[39][36] = 8'd155;
	sample_rom[39][37] = 8'd160;
	sample_rom[39][38] = 8'd156;
	sample_rom[39][39] = 8'd147;
	sample_rom[39][40] = 8'd133;
	sample_rom[39][41] = 8'd120;
	sample_rom[39][42] = 8'd108;
	sample_rom[39][43] = 8'd104;
	sample_rom[39][44] = 8'd109;
	sample_rom[39][45] = 8'd120;
	sample_rom[39][46] = 8'd135;
	sample_rom[39][47] = 8'd156;
	sample_rom[39][48] = 8'd173;
	sample_rom[39][49] = 8'd183;
	sample_rom[39][50] = 8'd187;
	sample_rom[39][51] = 8'd185;
	sample_rom[39][52] = 8'd174;
	sample_rom[39][53] = 8'd160;
	sample_rom[39][54] = 8'd142;
	sample_rom[39][55] = 8'd126;
	sample_rom[39][56] = 8'd115;
	sample_rom[39][57] = 8'd109;
	sample_rom[39][58] = 8'd105;
	sample_rom[39][59] = 8'd107;
	sample_rom[39][60] = 8'd110;
	sample_rom[39][61] = 8'd114;
	sample_rom[39][62] = 8'd118;
	sample_rom[39][63] = 8'd124;
	sample_rom[40][0] = 8'd131;
	sample_rom[40][1] = 8'd163;
	sample_rom[40][2] = 8'd194;
	sample_rom[40][3] = 8'd218;
	sample_rom[40][4] = 8'd233;
	sample_rom[40][5] = 8'd244;
	sample_rom[40][6] = 8'd245;
	sample_rom[40][7] = 8'd237;
	sample_rom[40][8] = 8'd224;
	sample_rom[40][9] = 8'd206;
	sample_rom[40][10] = 8'd185;
	sample_rom[40][11] = 8'd164;
	sample_rom[40][12] = 8'd144;
	sample_rom[40][13] = 8'd126;
	sample_rom[40][14] = 8'd113;
	sample_rom[40][15] = 8'd106;
	sample_rom[40][16] = 8'd103;
	sample_rom[40][17] = 8'd107;
	sample_rom[40][18] = 8'd112;
	sample_rom[40][19] = 8'd121;
	sample_rom[40][20] = 8'd133;
	sample_rom[40][21] = 8'd144;
	sample_rom[40][22] = 8'd154;
	sample_rom[40][23] = 8'd161;
	sample_rom[40][24] = 8'd166;
	sample_rom[40][25] = 8'd168;
	sample_rom[40][26] = 8'd169;
	sample_rom[40][27] = 8'd167;
	sample_rom[40][28] = 8'd163;
	sample_rom[40][29] = 8'd162;
	sample_rom[40][30] = 8'd158;
	sample_rom[40][31] = 8'd158;
	sample_rom[40][32] = 8'd156;
	sample_rom[40][33] = 8'd160;
	sample_rom[40][34] = 8'd161;
	sample_rom[40][35] = 8'd165;
	sample_rom[40][36] = 8'd168;
	sample_rom[40][37] = 8'd171;
	sample_rom[40][38] = 8'd172;
	sample_rom[40][39] = 8'd168;
	sample_rom[40][40] = 8'd166;
	sample_rom[40][41] = 8'd160;
	sample_rom[40][42] = 8'd154;
	sample_rom[40][43] = 8'd141;
	sample_rom[40][44] = 8'd132;
	sample_rom[40][45] = 8'd121;
	sample_rom[40][46] = 8'd111;
	sample_rom[40][47] = 8'd106;
	sample_rom[40][48] = 8'd102;
	sample_rom[40][49] = 8'd102;
	sample_rom[40][50] = 8'd108;
	sample_rom[40][51] = 8'd118;
	sample_rom[40][52] = 8'd130;
	sample_rom[40][53] = 8'd143;
	sample_rom[40][54] = 8'd157;
	sample_rom[40][55] = 8'd169;
	sample_rom[40][56] = 8'd181;
	sample_rom[40][57] = 8'd190;
	sample_rom[40][58] = 8'd194;
	sample_rom[40][59] = 8'd193;
	sample_rom[40][60] = 8'd187;
	sample_rom[40][61] = 8'd177;
	sample_rom[40][62] = 8'd161;
	sample_rom[40][63] = 8'd146;
	sample_rom[41][0] = 8'd130;
	sample_rom[41][1] = 8'd150;
	sample_rom[41][2] = 8'd166;
	sample_rom[41][3] = 8'd183;
	sample_rom[41][4] = 8'd196;
	sample_rom[41][5] = 8'd206;
	sample_rom[41][6] = 8'd211;
	sample_rom[41][7] = 8'd212;
	sample_rom[41][8] = 8'd211;
	sample_rom[41][9] = 8'd207;
	sample_rom[41][10] = 8'd201;
	sample_rom[41][11] = 8'd190;
	sample_rom[41][12] = 8'd181;
	sample_rom[41][13] = 8'd169;
	sample_rom[41][14] = 8'd158;
	sample_rom[41][15] = 8'd148;
	sample_rom[41][16] = 8'd140;
	sample_rom[41][17] = 8'd132;
	sample_rom[41][18] = 8'd126;
	sample_rom[41][19] = 8'd121;
	sample_rom[41][20] = 8'd118;
	sample_rom[41][21] = 8'd118;
	sample_rom[41][22] = 8'd116;
	sample_rom[41][23] = 8'd120;
	sample_rom[41][24] = 8'd120;
	sample_rom[41][25] = 8'd121;
	sample_rom[41][26] = 8'd124;
	sample_rom[41][27] = 8'd126;
	sample_rom[41][28] = 8'd127;
	sample_rom[41][29] = 8'd129;
	sample_rom[41][30] = 8'd129;
	sample_rom[41][31] = 8'd130;
	sample_rom[41][32] = 8'd130;
	sample_rom[41][33] = 8'd130;
	sample_rom[41][34] = 8'd129;
	sample_rom[41][35] = 8'd129;
	sample_rom[41][36] = 8'd128;
	sample_rom[41][37] = 8'd125;
	sample_rom[41][38] = 8'd124;
	sample_rom[41][39] = 8'd121;
	sample_rom[41][40] = 8'd120;
	sample_rom[41][41] = 8'd118;
	sample_rom[41][42] = 8'd119;
	sample_rom[41][43] = 8'd118;
	sample_rom[41][44] = 8'd120;
	sample_rom[41][45] = 8'd123;
	sample_rom[41][46] = 8'd127;
	sample_rom[41][47] = 8'd134;
	sample_rom[41][48] = 8'd140;
	sample_rom[41][49] = 8'd150;
	sample_rom[41][50] = 8'd160;
	sample_rom[41][51] = 8'd171;
	sample_rom[41][52] = 8'd181;
	sample_rom[41][53] = 8'd192;
	sample_rom[41][54] = 8'd201;
	sample_rom[41][55] = 8'd207;
	sample_rom[41][56] = 8'd210;
	sample_rom[41][57] = 8'd210;
	sample_rom[41][58] = 8'd209;
	sample_rom[41][59] = 8'd202;
	sample_rom[41][60] = 8'd192;
	sample_rom[41][61] = 8'd177;
	sample_rom[41][62] = 8'd161;
	sample_rom[41][63] = 8'd144;
	sample_rom[42][0] = 8'd130;
	sample_rom[42][1] = 8'd143;
	sample_rom[42][2] = 8'd154;
	sample_rom[42][3] = 8'd165;
	sample_rom[42][4] = 8'd175;
	sample_rom[42][5] = 8'd185;
	sample_rom[42][6] = 8'd195;
	sample_rom[42][7] = 8'd203;
	sample_rom[42][8] = 8'd210;
	sample_rom[42][9] = 8'd217;
	sample_rom[42][10] = 8'd221;
	sample_rom[42][11] = 8'd225;
	sample_rom[42][12] = 8'd227;
	sample_rom[42][13] = 8'd231;
	sample_rom[42][14] = 8'd230;
	sample_rom[42][15] = 8'd231;
	sample_rom[42][16] = 8'd229;
	sample_rom[42][17] = 8'd226;
	sample_rom[42][18] = 8'd223;
	sample_rom[42][19] = 8'd220;
	sample_rom[42][20] = 8'd215;
	sample_rom[42][21] = 8'd209;
	sample_rom[42][22] = 8'd203;
	sample_rom[42][23] = 8'd197;
	sample_rom[42][24] = 8'd190;
	sample_rom[42][25] = 8'd183;
	sample_rom[42][26] = 8'd176;
	sample_rom[42][27] = 8'd169;
	sample_rom[42][28] = 8'd163;
	sample_rom[42][29] = 8'd157;
	sample_rom[42][30] = 8'd152;
	sample_rom[42][31] = 8'd144;
	sample_rom[42][32] = 8'd140;
	sample_rom[42][33] = 8'd134;
	sample_rom[42][34] = 8'd129;
	sample_rom[42][35] = 8'd125;
	sample_rom[42][36] = 8'd121;
	sample_rom[42][37] = 8'd119;
	sample_rom[42][38] = 8'd115;
	sample_rom[42][39] = 8'd111;
	sample_rom[42][40] = 8'd110;
	sample_rom[42][41] = 8'd108;
	sample_rom[42][42] = 8'd108;
	sample_rom[42][43] = 8'd107;
	sample_rom[42][44] = 8'd107;
	sample_rom[42][45] = 8'd107;
	sample_rom[42][46] = 8'd105;
	sample_rom[42][47] = 8'd106;
	sample_rom[42][48] = 8'd106;
	sample_rom[42][49] = 8'd106;
	sample_rom[42][50] = 8'd109;
	sample_rom[42][51] = 8'd108;
	sample_rom[42][52] = 8'd110;
	sample_rom[42][53] = 8'd110;
	sample_rom[42][54] = 8'd112;
	sample_rom[42][55] = 8'd114;
	sample_rom[42][56] = 8'd115;
	sample_rom[42][57] = 8'd117;
	sample_rom[42][58] = 8'd118;
	sample_rom[42][59] = 8'd121;
	sample_rom[42][60] = 8'd121;
	sample_rom[42][61] = 8'd123;
	sample_rom[42][62] = 8'd124;
	sample_rom[42][63] = 8'd127;
	sample_rom[43][0] = 8'd131;
	sample_rom[43][1] = 8'd155;
	sample_rom[43][2] = 8'd179;
	sample_rom[43][3] = 8'd199;
	sample_rom[43][4] = 8'd214;
	sample_rom[43][5] = 8'd225;
	sample_rom[43][6] = 8'd233;
	sample_rom[43][7] = 8'd238;
	sample_rom[43][8] = 8'd234;
	sample_rom[43][9] = 8'd231;
	sample_rom[43][10] = 8'd225;
	sample_rom[43][11] = 8'd215;
	sample_rom[43][12] = 8'd206;
	sample_rom[43][13] = 8'd197;
	sample_rom[43][14] = 8'd189;
	sample_rom[43][15] = 8'd182;
	sample_rom[43][16] = 8'd174;
	sample_rom[43][17] = 8'd169;
	sample_rom[43][18] = 8'd165;
	sample_rom[43][19] = 8'd162;
	sample_rom[43][20] = 8'd158;
	sample_rom[43][21] = 8'd157;
	sample_rom[43][22] = 8'd153;
	sample_rom[43][23] = 8'd147;
	sample_rom[43][24] = 8'd140;
	sample_rom[43][25] = 8'd134;
	sample_rom[43][26] = 8'd127;
	sample_rom[43][27] = 8'd120;
	sample_rom[43][28] = 8'd113;
	sample_rom[43][29] = 8'd107;
	sample_rom[43][30] = 8'd103;
	sample_rom[43][31] = 8'd98;
	sample_rom[43][32] = 8'd99;
	sample_rom[43][33] = 8'd103;
	sample_rom[43][34] = 8'd106;
	sample_rom[43][35] = 8'd112;
	sample_rom[43][36] = 8'd118;
	sample_rom[43][37] = 8'd126;
	sample_rom[43][38] = 8'd132;
	sample_rom[43][39] = 8'd139;
	sample_rom[43][40] = 8'd144;
	sample_rom[43][41] = 8'd146;
	sample_rom[43][42] = 8'd147;
	sample_rom[43][43] = 8'd143;
	sample_rom[43][44] = 8'd140;
	sample_rom[43][45] = 8'd135;
	sample_rom[43][46] = 8'd127;
	sample_rom[43][47] = 8'd122;
	sample_rom[43][48] = 8'd114;
	sample_rom[43][49] = 8'd111;
	sample_rom[43][50] = 8'd107;
	sample_rom[43][51] = 8'd107;
	sample_rom[43][52] = 8'd107;
	sample_rom[43][53] = 8'd110;
	sample_rom[43][54] = 8'd114;
	sample_rom[43][55] = 8'd119;
	sample_rom[43][56] = 8'd124;
	sample_rom[43][57] = 8'd128;
	sample_rom[43][58] = 8'd131;
	sample_rom[43][59] = 8'd136;
	sample_rom[43][60] = 8'd136;
	sample_rom[43][61] = 8'd136;
	sample_rom[43][62] = 8'd134;
	sample_rom[43][63] = 8'd132;
	sample_rom[44][0] = 8'd130;
	sample_rom[44][1] = 8'd157;
	sample_rom[44][2] = 8'd180;
	sample_rom[44][3] = 8'd201;
	sample_rom[44][4] = 8'd217;
	sample_rom[44][5] = 8'd231;
	sample_rom[44][6] = 8'd238;
	sample_rom[44][7] = 8'd243;
	sample_rom[44][8] = 8'd241;
	sample_rom[44][9] = 8'd233;
	sample_rom[44][10] = 8'd224;
	sample_rom[44][11] = 8'd212;
	sample_rom[44][12] = 8'd194;
	sample_rom[44][13] = 8'd178;
	sample_rom[44][14] = 8'd161;
	sample_rom[44][15] = 8'd147;
	sample_rom[44][16] = 8'd131;
	sample_rom[44][17] = 8'd118;
	sample_rom[44][18] = 8'd108;
	sample_rom[44][19] = 8'd104;
	sample_rom[44][20] = 8'd101;
	sample_rom[44][21] = 8'd101;
	sample_rom[44][22] = 8'd104;
	sample_rom[44][23] = 8'd110;
	sample_rom[44][24] = 8'd116;
	sample_rom[44][25] = 8'd125;
	sample_rom[44][26] = 8'd134;
	sample_rom[44][27] = 8'd141;
	sample_rom[44][28] = 8'd146;
	sample_rom[44][29] = 8'd153;
	sample_rom[44][30] = 8'd155;
	sample_rom[44][31] = 8'd156;
	sample_rom[44][32] = 8'd157;
	sample_rom[44][33] = 8'd154;
	sample_rom[44][34] = 8'd150;
	sample_rom[44][35] = 8'd146;
	sample_rom[44][36] = 8'd142;
	sample_rom[44][37] = 8'd137;
	sample_rom[44][38] = 8'd130;
	sample_rom[44][39] = 8'd126;
	sample_rom[44][40] = 8'd123;
	sample_rom[44][41] = 8'd121;
	sample_rom[44][42] = 8'd119;
	sample_rom[44][43] = 8'd117;
	sample_rom[44][44] = 8'd118;
	sample_rom[44][45] = 8'd119;
	sample_rom[44][46] = 8'd119;
	sample_rom[44][47] = 8'd123;
	sample_rom[44][48] = 8'd125;
	sample_rom[44][49] = 8'd125;
	sample_rom[44][50] = 8'd129;
	sample_rom[44][51] = 8'd128;
	sample_rom[44][52] = 8'd130;
	sample_rom[44][53] = 8'd130;
	sample_rom[44][54] = 8'd129;
	sample_rom[44][55] = 8'd128;
	sample_rom[44][56] = 8'd128;
	sample_rom[44][57] = 8'd128;
	sample_rom[44][58] = 8'd128;
	sample_rom[44][59] = 8'd127;
	sample_rom[44][60] = 8'd126;
	sample_rom[44][61] = 8'd127;
	sample_rom[44][62] = 8'd127;
	sample_rom[44][63] = 8'd129;
	sample_rom[45][0] = 8'd131;
	sample_rom[45][1] = 8'd179;
	sample_rom[45][2] = 8'd217;
	sample_rom[45][3] = 8'd240;
	sample_rom[45][4] = 8'd244;
	sample_rom[45][5] = 8'd232;
	sample_rom[45][6] = 8'd208;
	sample_rom[45][7] = 8'd176;
	sample_rom[45][8] = 8'd150;
	sample_rom[45][9] = 8'd130;
	sample_rom[45][10] = 8'd125;
	sample_rom[45][11] = 8'd132;
	sample_rom[45][12] = 8'd154;
	sample_rom[45][13] = 8'd178;
	sample_rom[45][14] = 8'd206;
	sample_rom[45][15] = 8'd222;
	sample_rom[45][16] = 8'd227;
	sample_rom[45][17] = 8'd218;
	sample_rom[45][18] = 8'd193;
	sample_rom[45][19] = 8'd161;
	sample_rom[45][20] = 8'd128;
	sample_rom[45][21] = 8'd97;
	sample_rom[45][22] = 8'd77;
	sample_rom[45][23] = 8'd70;
	sample_rom[45][24] = 8'd76;
	sample_rom[45][25] = 8'd92;
	sample_rom[45][26] = 8'd116;
	sample_rom[45][27] = 8'd141;
	sample_rom[45][28] = 8'd160;
	sample_rom[45][29] = 8'd172;
	sample_rom[45][30] = 8'd173;
	sample_rom[45][31] = 8'd167;
	sample_rom[45][32] = 8'd155;
	sample_rom[45][33] = 8'd139;
	sample_rom[45][34] = 8'd124;
	sample_rom[45][35] = 8'd112;
	sample_rom[45][36] = 8'd108;
	sample_rom[45][37] = 8'd109;
	sample_rom[45][38] = 8'd114;
	sample_rom[45][39] = 8'd126;
	sample_rom[45][40] = 8'd135;
	sample_rom[45][41] = 8'd143;
	sample_rom[45][42] = 8'd150;
	sample_rom[45][43] = 8'd151;
	sample_rom[45][44] = 8'd149;
	sample_rom[45][45] = 8'd142;
	sample_rom[45][46] = 8'd133;
	sample_rom[45][47] = 8'd126;
	sample_rom[45][48] = 8'd121;
	sample_rom[45][49] = 8'd115;
	sample_rom[45][50] = 8'd115;
	sample_rom[45][51] = 8'd114;
	sample_rom[45][52] = 8'd118;
	sample_rom[45][53] = 8'd123;
	sample_rom[45][54] = 8'd127;
	sample_rom[45][55] = 8'd129;
	sample_rom[45][56] = 8'd135;
	sample_rom[45][57] = 8'd138;
	sample_rom[45][58] = 8'd139;
	sample_rom[45][59] = 8'd140;
	sample_rom[45][60] = 8'd140;
	sample_rom[45][61] = 8'd137;
	sample_rom[45][62] = 8'd136;
	sample_rom[45][63] = 8'd133;
	sample_rom[46][0] = 8'd130;
	sample_rom[46][1] = 8'd198;
	sample_rom[46][2] = 8'd236;
	sample_rom[46][3] = 8'd227;
	sample_rom[46][4] = 8'd182;
	sample_rom[46][5] = 8'd118;
	sample_rom[46][6] = 8'd68;
	sample_rom[46][7] = 8'd56;
	sample_rom[46][8] = 8'd84;
	sample_rom[46][9] = 8'd137;
	sample_rom[46][10] = 8'd195;
	sample_rom[46][11] = 8'd227;
	sample_rom[46][12] = 8'd227;
	sample_rom[46][13] = 8'd193;
	sample_rom[46][14] = 8'd150;
	sample_rom[46][15] = 8'd108;
	sample_rom[46][16] = 8'd86;
	sample_rom[46][17] = 8'd92;
	sample_rom[46][18] = 8'd114;
	sample_rom[46][19] = 8'd148;
	sample_rom[46][20] = 8'd172;
	sample_rom[46][21] = 8'd184;
	sample_rom[46][22] = 8'd171;
	sample_rom[46][23] = 8'd150;
	sample_rom[46][24] = 8'd122;
	sample_rom[46][25] = 8'd99;
	sample_rom[46][26] = 8'd89;
	sample_rom[46][27] = 8'd92;
	sample_rom[46][28] = 8'd106;
	sample_rom[46][29] = 8'd127;
	sample_rom[46][30] = 8'd142;
	sample_rom[46][31] = 8'd150;
	sample_rom[46][32] = 8'd144;
	sample_rom[46][33] = 8'd129;
	sample_rom[46][34] = 8'd110;
	sample_rom[46][35] = 8'd100;
	sample_rom[46][36] = 8'd97;
	sample_rom[46][37] = 8'd103;
	sample_rom[46][38] = 8'd119;
	sample_rom[46][39] = 8'd132;
	sample_rom[46][40] = 8'd140;
	sample_rom[46][41] = 8'd140;
	sample_rom[46][42] = 8'd135;
	sample_rom[46][43] = 8'd126;
	sample_rom[46][44] = 8'd122;
	sample_rom[46][45] = 8'd123;
	sample_rom[46][46] = 8'd127;
	sample_rom[46][47] = 8'd131;
	sample_rom[46][48] = 8'd135;
	sample_rom[46][49] = 8'd137;
	sample_rom[46][50] = 8'd137;
	sample_rom[46][51] = 8'd133;
	sample_rom[46][52] = 8'd133;
	sample_rom[46][53] = 8'd136;
	sample_rom[46][54] = 8'd135;
	sample_rom[46][55] = 8'd135;
	sample_rom[46][56] = 8'd133;
	sample_rom[46][57] = 8'd129;
	sample_rom[46][58] = 8'd128;
	sample_rom[46][59] = 8'd130;
	sample_rom[46][60] = 8'd131;
	sample_rom[46][61] = 8'd133;
	sample_rom[46][62] = 8'd135;
	sample_rom[46][63] = 8'd132;
	sample_rom[47][0] = 8'd131;
	sample_rom[47][1] = 8'd158;
	sample_rom[47][2] = 8'd178;
	sample_rom[47][3] = 8'd193;
	sample_rom[47][4] = 8'd195;
	sample_rom[47][5] = 8'd188;
	sample_rom[47][6] = 8'd177;
	sample_rom[47][7] = 8'd166;
	sample_rom[47][8] = 8'd160;
	sample_rom[47][9] = 8'd157;
	sample_rom[47][10] = 8'd163;
	sample_rom[47][11] = 8'd173;
	sample_rom[47][12] = 8'd185;
	sample_rom[47][13] = 8'd194;
	sample_rom[47][14] = 8'd196;
	sample_rom[47][15] = 8'd188;
	sample_rom[47][16] = 8'd171;
	sample_rom[47][17] = 8'd148;
	sample_rom[47][18] = 8'd124;
	sample_rom[47][19] = 8'd103;
	sample_rom[47][20] = 8'd90;
	sample_rom[47][21] = 8'd88;
	sample_rom[47][22] = 8'd93;
	sample_rom[47][23] = 8'd106;
	sample_rom[47][24] = 8'd122;
	sample_rom[47][25] = 8'd138;
	sample_rom[47][26] = 8'd147;
	sample_rom[47][27] = 8'd148;
	sample_rom[47][28] = 8'd143;
	sample_rom[47][29] = 8'd136;
	sample_rom[47][30] = 8'd127;
	sample_rom[47][31] = 8'd124;
	sample_rom[47][32] = 8'd129;
	sample_rom[47][33] = 8'd144;
	sample_rom[47][34] = 8'd164;
	sample_rom[47][35] = 8'd188;
	sample_rom[47][36] = 8'd211;
	sample_rom[47][37] = 8'd226;
	sample_rom[47][38] = 8'd232;
	sample_rom[47][39] = 8'd227;
	sample_rom[47][40] = 8'd216;
	sample_rom[47][41] = 8'd195;
	sample_rom[47][42] = 8'd178;
	sample_rom[47][43] = 8'd163;
	sample_rom[47][44] = 8'd156;
	sample_rom[47][45] = 8'd155;
	sample_rom[47][46] = 8'd160;
	sample_rom[47][47] = 8'd166;
	sample_rom[47][48] = 8'd171;
	sample_rom[47][49] = 8'd168;
	sample_rom[47][50] = 8'd159;
	sample_rom[47][51] = 8'd140;
	sample_rom[47][52] = 8'd116;
	sample_rom[47][53] = 8'd93;
	sample_rom[47][54] = 8'd74;
	sample_rom[47][55] = 8'd63;
	sample_rom[47][56] = 8'd64;
	sample_rom[47][57] = 8'd75;
	sample_rom[47][58] = 8'd91;
	sample_rom[47][59] = 8'd110;
	sample_rom[47][60] = 8'd128;
	sample_rom[47][61] = 8'd139;
	sample_rom[47][62] = 8'd141;
	sample_rom[47][63] = 8'd137;
	sample_rom[48][0] = 8'd131;
	sample_rom[48][1] = 8'd219;
	sample_rom[48][2] = 8'd238;
	sample_rom[48][3] = 8'd215;
	sample_rom[48][4] = 8'd208;
	sample_rom[48][5] = 8'd220;
	sample_rom[48][6] = 8'd210;
	sample_rom[48][7] = 8'd188;
	sample_rom[48][8] = 8'd185;
	sample_rom[48][9] = 8'd192;
	sample_rom[48][10] = 8'd190;
	sample_rom[48][11] = 8'd179;
	sample_rom[48][12] = 8'd178;
	sample_rom[48][13] = 8'd177;
	sample_rom[48][14] = 8'd166;
	sample_rom[48][15] = 8'd154;
	sample_rom[48][16] = 8'd157;
	sample_rom[48][17] = 8'd161;
	sample_rom[48][18] = 8'd158;
	sample_rom[48][19] = 8'd153;
	sample_rom[48][20] = 8'd157;
	sample_rom[48][21] = 8'd156;
	sample_rom[48][22] = 8'd140;
	sample_rom[48][23] = 8'd133;
	sample_rom[48][24] = 8'd140;
	sample_rom[48][25] = 8'd141;
	sample_rom[48][26] = 8'd133;
	sample_rom[48][27] = 8'd140;
	sample_rom[48][28] = 8'd162;
	sample_rom[48][29] = 8'd155;
	sample_rom[48][30] = 8'd113;
	sample_rom[48][31] = 8'd103;
	sample_rom[48][32] = 8'd148;
	sample_rom[48][33] = 8'd190;
	sample_rom[48][34] = 8'd177;
	sample_rom[48][35] = 8'd136;
	sample_rom[48][36] = 8'd129;
	sample_rom[48][37] = 8'd148;
	sample_rom[48][38] = 8'd150;
	sample_rom[48][39] = 8'd140;
	sample_rom[48][40] = 8'd137;
	sample_rom[48][41] = 8'd143;
	sample_rom[48][42] = 8'd134;
	sample_rom[48][43] = 8'd122;
	sample_rom[48][44] = 8'd121;
	sample_rom[48][45] = 8'd128;
	sample_rom[48][46] = 8'd128;
	sample_rom[48][47] = 8'd128;
	sample_rom[48][48] = 8'd136;
	sample_rom[48][49] = 8'd145;
	sample_rom[48][50] = 8'd141;
	sample_rom[48][51] = 8'd132;
	sample_rom[48][52] = 8'd137;
	sample_rom[48][53] = 8'd139;
	sample_rom[48][54] = 8'd131;
	sample_rom[48][55] = 8'd129;
	sample_rom[48][56] = 8'd138;
	sample_rom[48][57] = 8'd129;
	sample_rom[48][58] = 8'd104;
	sample_rom[48][59] = 8'd91;
	sample_rom[48][60] = 8'd94;
	sample_rom[48][61] = 8'd79;
	sample_rom[48][62] = 8'd47;
	sample_rom[48][63] = 8'd57;
	sample_rom[49][0] = 8'd133;
	sample_rom[49][1] = 8'd190;
	sample_rom[49][2] = 8'd206;
	sample_rom[49][3] = 8'd203;
	sample_rom[49][4] = 8'd213;
	sample_rom[49][5] = 8'd218;
	sample_rom[49][6] = 8'd197;
	sample_rom[49][7] = 8'd183;
	sample_rom[49][8] = 8'd205;
	sample_rom[49][9] = 8'd224;
	sample_rom[49][10] = 8'd205;
	sample_rom[49][11] = 8'd175;
	sample_rom[49][12] = 8'd170;
	sample_rom[49][13] = 8'd170;
	sample_rom[49][14] = 8'd153;
	sample_rom[49][15] = 8'd154;
	sample_rom[49][16] = 8'd194;
	sample_rom[49][17] = 8'd232;
	sample_rom[49][18] = 8'd231;
	sample_rom[49][19] = 8'd212;
	sample_rom[49][20] = 8'd206;
	sample_rom[49][21] = 8'd197;
	sample_rom[49][22] = 8'd164;
	sample_rom[49][23] = 8'd141;
	sample_rom[49][24] = 8'd156;
	sample_rom[49][25] = 8'd171;
	sample_rom[49][26] = 8'd150;
	sample_rom[49][27] = 8'd120;
	sample_rom[49][28] = 8'd117;
	sample_rom[49][29] = 8'd120;
	sample_rom[49][30] = 8'd111;
	sample_rom[49][31] = 8'd118;
	sample_rom[49][32] = 8'd167;
	sample_rom[49][33] = 8'd215;
	sample_rom[49][34] = 8'd221;
	sample_rom[49][35] = 8'd210;
	sample_rom[49][36] = 8'd212;
	sample_rom[49][37] = 8'd207;
	sample_rom[49][38] = 8'd178;
	sample_rom[49][39] = 8'd156;
	sample_rom[49][40] = 8'd169;
	sample_rom[49][41] = 8'd182;
	sample_rom[49][42] = 8'd156;
	sample_rom[49][43] = 8'd119;
	sample_rom[49][44] = 8'd108;
	sample_rom[49][45] = 8'd103;
	sample_rom[49][46] = 8'd82;
	sample_rom[49][47] = 8'd80;
	sample_rom[49][48] = 8'd118;
	sample_rom[49][49] = 8'd154;
	sample_rom[49][50] = 8'd152;
	sample_rom[49][51] = 8'd130;
	sample_rom[49][52] = 8'd126;
	sample_rom[49][53] = 8'd118;
	sample_rom[49][54] = 8'd87;
	sample_rom[49][55] = 8'd64;
	sample_rom[49][56] = 8'd81;
	sample_rom[49][57] = 8'd99;
	sample_rom[49][58] = 8'd82;
	sample_rom[49][59] = 8'd58;
	sample_rom[49][60] = 8'd59;
	sample_rom[49][61] = 8'd68;
	sample_rom[49][62] = 8'd63;
	sample_rom[49][63] = 8'd76;
	sample_rom[50][0] = 8'd128;
	sample_rom[50][1] = 8'd128;
	sample_rom[50][2] = 8'd128;
	sample_rom[50][3] = 8'd128;
	sample_rom[50][4] = 8'd128;
	sample_rom[50][5] = 8'd128;
	sample_rom[50][6] = 8'd128;
	sample_rom[50][7] = 8'd128;
	sample_rom[50][8] = 8'd128;
	sample_rom[50][9] = 8'd128;
	sample_rom[50][10] = 8'd128;
	sample_rom[50][11] = 8'd128;
	sample_rom[50][12] = 8'd128;
	sample_rom[50][13] = 8'd128;
	sample_rom[50][14] = 8'd128;
	sample_rom[50][15] = 8'd128;
	sample_rom[50][16] = 8'd128;
	sample_rom[50][17] = 8'd128;
	sample_rom[50][18] = 8'd128;
	sample_rom[50][19] = 8'd128;
	sample_rom[50][20] = 8'd128;
	sample_rom[50][21] = 8'd128;
	sample_rom[50][22] = 8'd128;
	sample_rom[50][23] = 8'd128;
	sample_rom[50][24] = 8'd128;
	sample_rom[50][25] = 8'd128;
	sample_rom[50][26] = 8'd128;
	sample_rom[50][27] = 8'd128;
	sample_rom[50][28] = 8'd128;
	sample_rom[50][29] = 8'd128;
	sample_rom[50][30] = 8'd128;
	sample_rom[50][31] = 8'd128;
	sample_rom[50][32] = 8'd128;
	sample_rom[50][33] = 8'd128;
	sample_rom[50][34] = 8'd128;
	sample_rom[50][35] = 8'd128;
	sample_rom[50][36] = 8'd128;
	sample_rom[50][37] = 8'd128;
	sample_rom[50][38] = 8'd128;
	sample_rom[50][39] = 8'd128;
	sample_rom[50][40] = 8'd128;
	sample_rom[50][41] = 8'd128;
	sample_rom[50][42] = 8'd128;
	sample_rom[50][43] = 8'd128;
	sample_rom[50][44] = 8'd128;
	sample_rom[50][45] = 8'd128;
	sample_rom[50][46] = 8'd128;
	sample_rom[50][47] = 8'd128;
	sample_rom[50][48] = 8'd128;
	sample_rom[50][49] = 8'd128;
	sample_rom[50][50] = 8'd128;
	sample_rom[50][51] = 8'd128;
	sample_rom[50][52] = 8'd128;
	sample_rom[50][53] = 8'd128;
	sample_rom[50][54] = 8'd128;
	sample_rom[50][55] = 8'd128;
	sample_rom[50][56] = 8'd128;
	sample_rom[50][57] = 8'd128;
	sample_rom[50][58] = 8'd128;
	sample_rom[50][59] = 8'd128;
	sample_rom[50][60] = 8'd128;
	sample_rom[50][61] = 8'd128;
	sample_rom[50][62] = 8'd128;
	sample_rom[50][63] = 8'd128;
	sample_rom[51][0] = 8'd128;
	sample_rom[51][1] = 8'd128;
	sample_rom[51][2] = 8'd128;
	sample_rom[51][3] = 8'd128;
	sample_rom[51][4] = 8'd128;
	sample_rom[51][5] = 8'd128;
	sample_rom[51][6] = 8'd128;
	sample_rom[51][7] = 8'd128;
	sample_rom[51][8] = 8'd128;
	sample_rom[51][9] = 8'd128;
	sample_rom[51][10] = 8'd128;
	sample_rom[51][11] = 8'd128;
	sample_rom[51][12] = 8'd128;
	sample_rom[51][13] = 8'd128;
	sample_rom[51][14] = 8'd128;
	sample_rom[51][15] = 8'd128;
	sample_rom[51][16] = 8'd128;
	sample_rom[51][17] = 8'd128;
	sample_rom[51][18] = 8'd128;
	sample_rom[51][19] = 8'd128;
	sample_rom[51][20] = 8'd128;
	sample_rom[51][21] = 8'd128;
	sample_rom[51][22] = 8'd128;
	sample_rom[51][23] = 8'd128;
	sample_rom[51][24] = 8'd128;
	sample_rom[51][25] = 8'd128;
	sample_rom[51][26] = 8'd128;
	sample_rom[51][27] = 8'd128;
	sample_rom[51][28] = 8'd128;
	sample_rom[51][29] = 8'd128;
	sample_rom[51][30] = 8'd128;
	sample_rom[51][31] = 8'd128;
	sample_rom[51][32] = 8'd128;
	sample_rom[51][33] = 8'd128;
	sample_rom[51][34] = 8'd128;
	sample_rom[51][35] = 8'd128;
	sample_rom[51][36] = 8'd128;
	sample_rom[51][37] = 8'd128;
	sample_rom[51][38] = 8'd128;
	sample_rom[51][39] = 8'd128;
	sample_rom[51][40] = 8'd128;
	sample_rom[51][41] = 8'd128;
	sample_rom[51][42] = 8'd128;
	sample_rom[51][43] = 8'd128;
	sample_rom[51][44] = 8'd128;
	sample_rom[51][45] = 8'd128;
	sample_rom[51][46] = 8'd128;
	sample_rom[51][47] = 8'd128;
	sample_rom[51][48] = 8'd128;
	sample_rom[51][49] = 8'd128;
	sample_rom[51][50] = 8'd128;
	sample_rom[51][51] = 8'd128;
	sample_rom[51][52] = 8'd128;
	sample_rom[51][53] = 8'd128;
	sample_rom[51][54] = 8'd128;
	sample_rom[51][55] = 8'd128;
	sample_rom[51][56] = 8'd128;
	sample_rom[51][57] = 8'd128;
	sample_rom[51][58] = 8'd128;
	sample_rom[51][59] = 8'd128;
	sample_rom[51][60] = 8'd128;
	sample_rom[51][61] = 8'd128;
	sample_rom[51][62] = 8'd128;
	sample_rom[51][63] = 8'd128;
	sample_rom[52][0] = 8'd128;
	sample_rom[52][1] = 8'd128;
	sample_rom[52][2] = 8'd128;
	sample_rom[52][3] = 8'd128;
	sample_rom[52][4] = 8'd128;
	sample_rom[52][5] = 8'd128;
	sample_rom[52][6] = 8'd128;
	sample_rom[52][7] = 8'd128;
	sample_rom[52][8] = 8'd128;
	sample_rom[52][9] = 8'd128;
	sample_rom[52][10] = 8'd128;
	sample_rom[52][11] = 8'd128;
	sample_rom[52][12] = 8'd128;
	sample_rom[52][13] = 8'd128;
	sample_rom[52][14] = 8'd128;
	sample_rom[52][15] = 8'd128;
	sample_rom[52][16] = 8'd128;
	sample_rom[52][17] = 8'd128;
	sample_rom[52][18] = 8'd128;
	sample_rom[52][19] = 8'd128;
	sample_rom[52][20] = 8'd128;
	sample_rom[52][21] = 8'd128;
	sample_rom[52][22] = 8'd128;
	sample_rom[52][23] = 8'd128;
	sample_rom[52][24] = 8'd128;
	sample_rom[52][25] = 8'd128;
	sample_rom[52][26] = 8'd128;
	sample_rom[52][27] = 8'd128;
	sample_rom[52][28] = 8'd128;
	sample_rom[52][29] = 8'd128;
	sample_rom[52][30] = 8'd128;
	sample_rom[52][31] = 8'd128;
	sample_rom[52][32] = 8'd128;
	sample_rom[52][33] = 8'd128;
	sample_rom[52][34] = 8'd128;
	sample_rom[52][35] = 8'd128;
	sample_rom[52][36] = 8'd128;
	sample_rom[52][37] = 8'd128;
	sample_rom[52][38] = 8'd128;
	sample_rom[52][39] = 8'd128;
	sample_rom[52][40] = 8'd128;
	sample_rom[52][41] = 8'd128;
	sample_rom[52][42] = 8'd128;
	sample_rom[52][43] = 8'd128;
	sample_rom[52][44] = 8'd128;
	sample_rom[52][45] = 8'd128;
	sample_rom[52][46] = 8'd128;
	sample_rom[52][47] = 8'd128;
	sample_rom[52][48] = 8'd128;
	sample_rom[52][49] = 8'd128;
	sample_rom[52][50] = 8'd128;
	sample_rom[52][51] = 8'd128;
	sample_rom[52][52] = 8'd128;
	sample_rom[52][53] = 8'd128;
	sample_rom[52][54] = 8'd128;
	sample_rom[52][55] = 8'd128;
	sample_rom[52][56] = 8'd128;
	sample_rom[52][57] = 8'd128;
	sample_rom[52][58] = 8'd128;
	sample_rom[52][59] = 8'd128;
	sample_rom[52][60] = 8'd128;
	sample_rom[52][61] = 8'd128;
	sample_rom[52][62] = 8'd128;
	sample_rom[52][63] = 8'd128;
	sample_rom[53][0] = 8'd130;
	sample_rom[53][1] = 8'd207;
	sample_rom[53][2] = 8'd241;
	sample_rom[53][3] = 8'd238;
	sample_rom[53][4] = 8'd222;
	sample_rom[53][5] = 8'd214;
	sample_rom[53][6] = 8'd218;
	sample_rom[53][7] = 8'd226;
	sample_rom[53][8] = 8'd223;
	sample_rom[53][9] = 8'd214;
	sample_rom[53][10] = 8'd211;
	sample_rom[53][11] = 8'd213;
	sample_rom[53][12] = 8'd214;
	sample_rom[53][13] = 8'd210;
	sample_rom[53][14] = 8'd203;
	sample_rom[53][15] = 8'd197;
	sample_rom[53][16] = 8'd198;
	sample_rom[53][17] = 8'd202;
	sample_rom[53][18] = 8'd203;
	sample_rom[53][19] = 8'd196;
	sample_rom[53][20] = 8'd192;
	sample_rom[53][21] = 8'd195;
	sample_rom[53][22] = 8'd195;
	sample_rom[53][23] = 8'd189;
	sample_rom[53][24] = 8'd186;
	sample_rom[53][25] = 8'd183;
	sample_rom[53][26] = 8'd184;
	sample_rom[53][27] = 8'd185;
	sample_rom[53][28] = 8'd187;
	sample_rom[53][29] = 8'd181;
	sample_rom[53][30] = 8'd180;
	sample_rom[53][31] = 8'd176;
	sample_rom[53][32] = 8'd178;
	sample_rom[53][33] = 8'd183;
	sample_rom[53][34] = 8'd176;
	sample_rom[53][35] = 8'd173;
	sample_rom[53][36] = 8'd175;
	sample_rom[53][37] = 8'd170;
	sample_rom[53][38] = 8'd169;
	sample_rom[53][39] = 8'd166;
	sample_rom[53][40] = 8'd163;
	sample_rom[53][41] = 8'd160;
	sample_rom[53][42] = 8'd163;
	sample_rom[53][43] = 8'd158;
	sample_rom[53][44] = 8'd157;
	sample_rom[53][45] = 8'd157;
	sample_rom[53][46] = 8'd151;
	sample_rom[53][47] = 8'd155;
	sample_rom[53][48] = 8'd153;
	sample_rom[53][49] = 8'd151;
	sample_rom[53][50] = 8'd150;
	sample_rom[53][51] = 8'd150;
	sample_rom[53][52] = 8'd152;
	sample_rom[53][53] = 8'd147;
	sample_rom[53][54] = 8'd141;
	sample_rom[53][55] = 8'd140;
	sample_rom[53][56] = 8'd137;
	sample_rom[53][57] = 8'd135;
	sample_rom[53][58] = 8'd135;
	sample_rom[53][59] = 8'd130;
	sample_rom[53][60] = 8'd124;
	sample_rom[53][61] = 8'd125;
	sample_rom[53][62] = 8'd126;
	sample_rom[53][63] = 8'd129;
	sample_rom[54][0] = 8'd131;
	sample_rom[54][1] = 8'd139;
	sample_rom[54][2] = 8'd147;
	sample_rom[54][3] = 8'd154;
	sample_rom[54][4] = 8'd160;
	sample_rom[54][5] = 8'd165;
	sample_rom[54][6] = 8'd173;
	sample_rom[54][7] = 8'd179;
	sample_rom[54][8] = 8'd185;
	sample_rom[54][9] = 8'd191;
	sample_rom[54][10] = 8'd197;
	sample_rom[54][11] = 8'd203;
	sample_rom[54][12] = 8'd207;
	sample_rom[54][13] = 8'd212;
	sample_rom[54][14] = 8'd216;
	sample_rom[54][15] = 8'd221;
	sample_rom[54][16] = 8'd223;
	sample_rom[54][17] = 8'd226;
	sample_rom[54][18] = 8'd226;
	sample_rom[54][19] = 8'd228;
	sample_rom[54][20] = 8'd229;
	sample_rom[54][21] = 8'd231;
	sample_rom[54][22] = 8'd231;
	sample_rom[54][23] = 8'd232;
	sample_rom[54][24] = 8'd232;
	sample_rom[54][25] = 8'd232;
	sample_rom[54][26] = 8'd230;
	sample_rom[54][27] = 8'd229;
	sample_rom[54][28] = 8'd227;
	sample_rom[54][29] = 8'd226;
	sample_rom[54][30] = 8'd223;
	sample_rom[54][31] = 8'd221;
	sample_rom[54][32] = 8'd218;
	sample_rom[54][33] = 8'd215;
	sample_rom[54][34] = 8'd212;
	sample_rom[54][35] = 8'd209;
	sample_rom[54][36] = 8'd206;
	sample_rom[54][37] = 8'd202;
	sample_rom[54][38] = 8'd198;
	sample_rom[54][39] = 8'd194;
	sample_rom[54][40] = 8'd190;
	sample_rom[54][41] = 8'd187;
	sample_rom[54][42] = 8'd183;
	sample_rom[54][43] = 8'd178;
	sample_rom[54][44] = 8'd175;
	sample_rom[54][45] = 8'd171;
	sample_rom[54][46] = 8'd170;
	sample_rom[54][47] = 8'd166;
	sample_rom[54][48] = 8'd163;
	sample_rom[54][49] = 8'd160;
	sample_rom[54][50] = 8'd157;
	sample_rom[54][51] = 8'd154;
	sample_rom[54][52] = 8'd152;
	sample_rom[54][53] = 8'd149;
	sample_rom[54][54] = 8'd146;
	sample_rom[54][55] = 8'd143;
	sample_rom[54][56] = 8'd141;
	sample_rom[54][57] = 8'd139;
	sample_rom[54][58] = 8'd137;
	sample_rom[54][59] = 8'd136;
	sample_rom[54][60] = 8'd135;
	sample_rom[54][61] = 8'd133;
	sample_rom[54][62] = 8'd130;
	sample_rom[54][63] = 8'd128;
	sample_rom[55][0] = 8'd131;
	sample_rom[55][1] = 8'd140;
	sample_rom[55][2] = 8'd150;
	sample_rom[55][3] = 8'd158;
	sample_rom[55][4] = 8'd166;
	sample_rom[55][5] = 8'd173;
	sample_rom[55][6] = 8'd182;
	sample_rom[55][7] = 8'd189;
	sample_rom[55][8] = 8'd195;
	sample_rom[55][9] = 8'd203;
	sample_rom[55][10] = 8'd209;
	sample_rom[55][11] = 8'd214;
	sample_rom[55][12] = 8'd220;
	sample_rom[55][13] = 8'd223;
	sample_rom[55][14] = 8'd228;
	sample_rom[55][15] = 8'd232;
	sample_rom[55][16] = 8'd234;
	sample_rom[55][17] = 8'd237;
	sample_rom[55][18] = 8'd238;
	sample_rom[55][19] = 8'd239;
	sample_rom[55][20] = 8'd238;
	sample_rom[55][21] = 8'd239;
	sample_rom[55][22] = 8'd239;
	sample_rom[55][23] = 8'd239;
	sample_rom[55][24] = 8'd236;
	sample_rom[55][25] = 8'd234;
	sample_rom[55][26] = 8'd232;
	sample_rom[55][27] = 8'd229;
	sample_rom[55][28] = 8'd225;
	sample_rom[55][29] = 8'd223;
	sample_rom[55][30] = 8'd219;
	sample_rom[55][31] = 8'd214;
	sample_rom[55][32] = 8'd210;
	sample_rom[55][33] = 8'd205;
	sample_rom[55][34] = 8'd201;
	sample_rom[55][35] = 8'd196;
	sample_rom[55][36] = 8'd191;
	sample_rom[55][37] = 8'd187;
	sample_rom[55][38] = 8'd182;
	sample_rom[55][39] = 8'd177;
	sample_rom[55][40] = 8'd173;
	sample_rom[55][41] = 8'd170;
	sample_rom[55][42] = 8'd165;
	sample_rom[55][43] = 8'd160;
	sample_rom[55][44] = 8'd157;
	sample_rom[55][45] = 8'd155;
	sample_rom[55][46] = 8'd152;
	sample_rom[55][47] = 8'd148;
	sample_rom[55][48] = 8'd145;
	sample_rom[55][49] = 8'd143;
	sample_rom[55][50] = 8'd140;
	sample_rom[55][51] = 8'd138;
	sample_rom[55][52] = 8'd136;
	sample_rom[55][53] = 8'd135;
	sample_rom[55][54] = 8'd133;
	sample_rom[55][55] = 8'd131;
	sample_rom[55][56] = 8'd130;
	sample_rom[55][57] = 8'd130;
	sample_rom[55][58] = 8'd128;
	sample_rom[55][59] = 8'd129;
	sample_rom[55][60] = 8'd128;
	sample_rom[55][61] = 8'd129;
	sample_rom[55][62] = 8'd127;
	sample_rom[55][63] = 8'd127;
	sample_rom[56][0] = 8'd131;
	sample_rom[56][1] = 8'd146;
	sample_rom[56][2] = 8'd159;
	sample_rom[56][3] = 8'd168;
	sample_rom[56][4] = 8'd180;
	sample_rom[56][5] = 8'd190;
	sample_rom[56][6] = 8'd201;
	sample_rom[56][7] = 8'd209;
	sample_rom[56][8] = 8'd218;
	sample_rom[56][9] = 8'd224;
	sample_rom[56][10] = 8'd231;
	sample_rom[56][11] = 8'd236;
	sample_rom[56][12] = 8'd240;
	sample_rom[56][13] = 8'd243;
	sample_rom[56][14] = 8'd245;
	sample_rom[56][15] = 8'd249;
	sample_rom[56][16] = 8'd250;
	sample_rom[56][17] = 8'd249;
	sample_rom[56][18] = 8'd246;
	sample_rom[56][19] = 8'd246;
	sample_rom[56][20] = 8'd243;
	sample_rom[56][21] = 8'd241;
	sample_rom[56][22] = 8'd239;
	sample_rom[56][23] = 8'd236;
	sample_rom[56][24] = 8'd233;
	sample_rom[56][25] = 8'd231;
	sample_rom[56][26] = 8'd227;
	sample_rom[56][27] = 8'd223;
	sample_rom[56][28] = 8'd220;
	sample_rom[56][29] = 8'd216;
	sample_rom[56][30] = 8'd213;
	sample_rom[56][31] = 8'd208;
	sample_rom[56][32] = 8'd205;
	sample_rom[56][33] = 8'd201;
	sample_rom[56][34] = 8'd198;
	sample_rom[56][35] = 8'd193;
	sample_rom[56][36] = 8'd191;
	sample_rom[56][37] = 8'd186;
	sample_rom[56][38] = 8'd183;
	sample_rom[56][39] = 8'd179;
	sample_rom[56][40] = 8'd175;
	sample_rom[56][41] = 8'd173;
	sample_rom[56][42] = 8'd170;
	sample_rom[56][43] = 8'd165;
	sample_rom[56][44] = 8'd164;
	sample_rom[56][45] = 8'd161;
	sample_rom[56][46] = 8'd160;
	sample_rom[56][47] = 8'd159;
	sample_rom[56][48] = 8'd157;
	sample_rom[56][49] = 8'd154;
	sample_rom[56][50] = 8'd152;
	sample_rom[56][51] = 8'd150;
	sample_rom[56][52] = 8'd148;
	sample_rom[56][53] = 8'd147;
	sample_rom[56][54] = 8'd144;
	sample_rom[56][55] = 8'd143;
	sample_rom[56][56] = 8'd141;
	sample_rom[56][57] = 8'd140;
	sample_rom[56][58] = 8'd138;
	sample_rom[56][59] = 8'd137;
	sample_rom[56][60] = 8'd136;
	sample_rom[56][61] = 8'd133;
	sample_rom[56][62] = 8'd131;
	sample_rom[56][63] = 8'd128;
	sample_rom[57][0] = 8'd132;
	sample_rom[57][1] = 8'd149;
	sample_rom[57][2] = 8'd165;
	sample_rom[57][3] = 8'd179;
	sample_rom[57][4] = 8'd194;
	sample_rom[57][5] = 8'd206;
	sample_rom[57][6] = 8'd217;
	sample_rom[57][7] = 8'd223;
	sample_rom[57][8] = 8'd232;
	sample_rom[57][9] = 8'd236;
	sample_rom[57][10] = 8'd239;
	sample_rom[57][11] = 8'd242;
	sample_rom[57][12] = 8'd241;
	sample_rom[57][13] = 8'd240;
	sample_rom[57][14] = 8'd238;
	sample_rom[57][15] = 8'd237;
	sample_rom[57][16] = 8'd235;
	sample_rom[57][17] = 8'd232;
	sample_rom[57][18] = 8'd227;
	sample_rom[57][19] = 8'd223;
	sample_rom[57][20] = 8'd221;
	sample_rom[57][21] = 8'd219;
	sample_rom[57][22] = 8'd215;
	sample_rom[57][23] = 8'd211;
	sample_rom[57][24] = 8'd208;
	sample_rom[57][25] = 8'd205;
	sample_rom[57][26] = 8'd202;
	sample_rom[57][27] = 8'd198;
	sample_rom[57][28] = 8'd196;
	sample_rom[57][29] = 8'd192;
	sample_rom[57][30] = 8'd189;
	sample_rom[57][31] = 8'd184;
	sample_rom[57][32] = 8'd182;
	sample_rom[57][33] = 8'd178;
	sample_rom[57][34] = 8'd174;
	sample_rom[57][35] = 8'd171;
	sample_rom[57][36] = 8'd168;
	sample_rom[57][37] = 8'd163;
	sample_rom[57][38] = 8'd160;
	sample_rom[57][39] = 8'd158;
	sample_rom[57][40] = 8'd154;
	sample_rom[57][41] = 8'd152;
	sample_rom[57][42] = 8'd149;
	sample_rom[57][43] = 8'd147;
	sample_rom[57][44] = 8'd144;
	sample_rom[57][45] = 8'd142;
	sample_rom[57][46] = 8'd143;
	sample_rom[57][47] = 8'd142;
	sample_rom[57][48] = 8'd144;
	sample_rom[57][49] = 8'd143;
	sample_rom[57][50] = 8'd145;
	sample_rom[57][51] = 8'd147;
	sample_rom[57][52] = 8'd148;
	sample_rom[57][53] = 8'd150;
	sample_rom[57][54] = 8'd154;
	sample_rom[57][55] = 8'd151;
	sample_rom[57][56] = 8'd153;
	sample_rom[57][57] = 8'd152;
	sample_rom[57][58] = 8'd151;
	sample_rom[57][59] = 8'd150;
	sample_rom[57][60] = 8'd146;
	sample_rom[57][61] = 8'd144;
	sample_rom[57][62] = 8'd136;
	sample_rom[57][63] = 8'd134;
	sample_rom[58][0] = 8'd130;
	sample_rom[58][1] = 8'd150;
	sample_rom[58][2] = 8'd166;
	sample_rom[58][3] = 8'd180;
	sample_rom[58][4] = 8'd190;
	sample_rom[58][5] = 8'd193;
	sample_rom[58][6] = 8'd195;
	sample_rom[58][7] = 8'd193;
	sample_rom[58][8] = 8'd192;
	sample_rom[58][9] = 8'd189;
	sample_rom[58][10] = 8'd187;
	sample_rom[58][11] = 8'd186;
	sample_rom[58][12] = 8'd182;
	sample_rom[58][13] = 8'd182;
	sample_rom[58][14] = 8'd184;
	sample_rom[58][15] = 8'd185;
	sample_rom[58][16] = 8'd184;
	sample_rom[58][17] = 8'd183;
	sample_rom[58][18] = 8'd182;
	sample_rom[58][19] = 8'd181;
	sample_rom[58][20] = 8'd181;
	sample_rom[58][21] = 8'd185;
	sample_rom[58][22] = 8'd188;
	sample_rom[58][23] = 8'd192;
	sample_rom[58][24] = 8'd200;
	sample_rom[58][25] = 8'd208;
	sample_rom[58][26] = 8'd215;
	sample_rom[58][27] = 8'd222;
	sample_rom[58][28] = 8'd229;
	sample_rom[58][29] = 8'd234;
	sample_rom[58][30] = 8'd234;
	sample_rom[58][31] = 8'd234;
	sample_rom[58][32] = 8'd234;
	sample_rom[58][33] = 8'd230;
	sample_rom[58][34] = 8'd227;
	sample_rom[58][35] = 8'd223;
	sample_rom[58][36] = 8'd219;
	sample_rom[58][37] = 8'd215;
	sample_rom[58][38] = 8'd213;
	sample_rom[58][39] = 8'd210;
	sample_rom[58][40] = 8'd207;
	sample_rom[58][41] = 8'd207;
	sample_rom[58][42] = 8'd206;
	sample_rom[58][43] = 8'd205;
	sample_rom[58][44] = 8'd205;
	sample_rom[58][45] = 8'd204;
	sample_rom[58][46] = 8'd205;
	sample_rom[58][47] = 8'd200;
	sample_rom[58][48] = 8'd197;
	sample_rom[58][49] = 8'd190;
	sample_rom[58][50] = 8'd183;
	sample_rom[58][51] = 8'd175;
	sample_rom[58][52] = 8'd168;
	sample_rom[58][53] = 8'd161;
	sample_rom[58][54] = 8'd156;
	sample_rom[58][55] = 8'd150;
	sample_rom[58][56] = 8'd147;
	sample_rom[58][57] = 8'd144;
	sample_rom[58][58] = 8'd142;
	sample_rom[58][59] = 8'd142;
	sample_rom[58][60] = 8'd140;
	sample_rom[58][61] = 8'd138;
	sample_rom[58][62] = 8'd133;
	sample_rom[58][63] = 8'd130;
	sample_rom[59][0] = 8'd131;
	sample_rom[59][1] = 8'd200;
	sample_rom[59][2] = 8'd236;
	sample_rom[59][3] = 8'd242;
	sample_rom[59][4] = 8'd221;
	sample_rom[59][5] = 8'd188;
	sample_rom[59][6] = 8'd160;
	sample_rom[59][7] = 8'd144;
	sample_rom[59][8] = 8'd144;
	sample_rom[59][9] = 8'd157;
	sample_rom[59][10] = 8'd168;
	sample_rom[59][11] = 8'd174;
	sample_rom[59][12] = 8'd177;
	sample_rom[59][13] = 8'd175;
	sample_rom[59][14] = 8'd179;
	sample_rom[59][15] = 8'd188;
	sample_rom[59][16] = 8'd202;
	sample_rom[59][17] = 8'd217;
	sample_rom[59][18] = 8'd225;
	sample_rom[59][19] = 8'd209;
	sample_rom[59][20] = 8'd179;
	sample_rom[59][21] = 8'd149;
	sample_rom[59][22] = 8'd121;
	sample_rom[59][23] = 8'd110;
	sample_rom[59][24] = 8'd116;
	sample_rom[59][25] = 8'd137;
	sample_rom[59][26] = 8'd166;
	sample_rom[59][27] = 8'd187;
	sample_rom[59][28] = 8'd192;
	sample_rom[59][29] = 8'd179;
	sample_rom[59][30] = 8'd160;
	sample_rom[59][31] = 8'd140;
	sample_rom[59][32] = 8'd129;
	sample_rom[59][33] = 8'd129;
	sample_rom[59][34] = 8'd142;
	sample_rom[59][35] = 8'd155;
	sample_rom[59][36] = 8'd160;
	sample_rom[59][37] = 8'd157;
	sample_rom[59][38] = 8'd144;
	sample_rom[59][39] = 8'd130;
	sample_rom[59][40] = 8'd123;
	sample_rom[59][41] = 8'd123;
	sample_rom[59][42] = 8'd136;
	sample_rom[59][43] = 8'd157;
	sample_rom[59][44] = 8'd170;
	sample_rom[59][45] = 8'd168;
	sample_rom[59][46] = 8'd159;
	sample_rom[59][47] = 8'd147;
	sample_rom[59][48] = 8'd138;
	sample_rom[59][49] = 8'd133;
	sample_rom[59][50] = 8'd136;
	sample_rom[59][51] = 8'd147;
	sample_rom[59][52] = 8'd156;
	sample_rom[59][53] = 8'd159;
	sample_rom[59][54] = 8'd148;
	sample_rom[59][55] = 8'd130;
	sample_rom[59][56] = 8'd117;
	sample_rom[59][57] = 8'd112;
	sample_rom[59][58] = 8'd113;
	sample_rom[59][59] = 8'd128;
	sample_rom[59][60] = 8'd143;
	sample_rom[59][61] = 8'd145;
	sample_rom[59][62] = 8'd145;
	sample_rom[59][63] = 8'd137;
	sample_rom[60][0] = 8'd130;
	sample_rom[60][1] = 8'd201;
	sample_rom[60][2] = 8'd236;
	sample_rom[60][3] = 8'd223;
	sample_rom[60][4] = 8'd168;
	sample_rom[60][5] = 8'd95;
	sample_rom[60][6] = 8'd38;
	sample_rom[60][7] = 8'd23;
	sample_rom[60][8] = 8'd55;
	sample_rom[60][9] = 8'd120;
	sample_rom[60][10] = 8'd188;
	sample_rom[60][11] = 8'd225;
	sample_rom[60][12] = 8'd219;
	sample_rom[60][13] = 8'd171;
	sample_rom[60][14] = 8'd107;
	sample_rom[60][15] = 8'd53;
	sample_rom[60][16] = 8'd33;
	sample_rom[60][17] = 8'd58;
	sample_rom[60][18] = 8'd111;
	sample_rom[60][19] = 8'd173;
	sample_rom[60][20] = 8'd211;
	sample_rom[60][21] = 8'd212;
	sample_rom[60][22] = 8'd173;
	sample_rom[60][23] = 8'd117;
	sample_rom[60][24] = 8'd68;
	sample_rom[60][25] = 8'd46;
	sample_rom[60][26] = 8'd63;
	sample_rom[60][27] = 8'd107;
	sample_rom[60][28] = 8'd160;
	sample_rom[60][29] = 8'd198;
	sample_rom[60][30] = 8'd204;
	sample_rom[60][31] = 8'd175;
	sample_rom[60][32] = 8'd126;
	sample_rom[60][33] = 8'd78;
	sample_rom[60][34] = 8'd55;
	sample_rom[60][35] = 8'd65;
	sample_rom[60][36] = 8'd102;
	sample_rom[60][37] = 8'd151;
	sample_rom[60][38] = 8'd186;
	sample_rom[60][39] = 8'd197;
	sample_rom[60][40] = 8'd176;
	sample_rom[60][41] = 8'd134;
	sample_rom[60][42] = 8'd91;
	sample_rom[60][43] = 8'd66;
	sample_rom[60][44] = 8'd71;
	sample_rom[60][45] = 8'd101;
	sample_rom[60][46] = 8'd143;
	sample_rom[60][47] = 8'd174;
	sample_rom[60][48] = 8'd184;
	sample_rom[60][49] = 8'd171;
	sample_rom[60][50] = 8'd139;
	sample_rom[60][51] = 8'd101;
	sample_rom[60][52] = 8'd81;
	sample_rom[60][53] = 8'd81;
	sample_rom[60][54] = 8'd102;
	sample_rom[60][55] = 8'd135;
	sample_rom[60][56] = 8'd162;
	sample_rom[60][57] = 8'd173;
	sample_rom[60][58] = 8'd164;
	sample_rom[60][59] = 8'd139;
	sample_rom[60][60] = 8'd112;
	sample_rom[60][61] = 8'd92;
	sample_rom[60][62] = 8'd88;
	sample_rom[60][63] = 8'd102;
	sample_rom[61][0] = 8'd131;
	sample_rom[61][1] = 8'd141;
	sample_rom[61][2] = 8'd149;
	sample_rom[61][3] = 8'd159;
	sample_rom[61][4] = 8'd166;
	sample_rom[61][5] = 8'd173;
	sample_rom[61][6] = 8'd181;
	sample_rom[61][7] = 8'd187;
	sample_rom[61][8] = 8'd193;
	sample_rom[61][9] = 8'd200;
	sample_rom[61][10] = 8'd205;
	sample_rom[61][11] = 8'd208;
	sample_rom[61][12] = 8'd212;
	sample_rom[61][13] = 8'd216;
	sample_rom[61][14] = 8'd218;
	sample_rom[61][15] = 8'd220;
	sample_rom[61][16] = 8'd221;
	sample_rom[61][17] = 8'd220;
	sample_rom[61][18] = 8'd220;
	sample_rom[61][19] = 8'd219;
	sample_rom[61][20] = 8'd217;
	sample_rom[61][21] = 8'd217;
	sample_rom[61][22] = 8'd214;
	sample_rom[61][23] = 8'd213;
	sample_rom[61][24] = 8'd210;
	sample_rom[61][25] = 8'd209;
	sample_rom[61][26] = 8'd206;
	sample_rom[61][27] = 8'd204;
	sample_rom[61][28] = 8'd203;
	sample_rom[61][29] = 8'd201;
	sample_rom[61][30] = 8'd201;
	sample_rom[61][31] = 8'd199;
	sample_rom[61][32] = 8'd199;
	sample_rom[61][33] = 8'd198;
	sample_rom[61][34] = 8'd198;
	sample_rom[61][35] = 8'd199;
	sample_rom[61][36] = 8'd198;
	sample_rom[61][37] = 8'd200;
	sample_rom[61][38] = 8'd200;
	sample_rom[61][39] = 8'd202;
	sample_rom[61][40] = 8'd204;
	sample_rom[61][41] = 8'd203;
	sample_rom[61][42] = 8'd206;
	sample_rom[61][43] = 8'd206;
	sample_rom[61][44] = 8'd208;
	sample_rom[61][45] = 8'd207;
	sample_rom[61][46] = 8'd208;
	sample_rom[61][47] = 8'd209;
	sample_rom[61][48] = 8'd209;
	sample_rom[61][49] = 8'd207;
	sample_rom[61][50] = 8'd205;
	sample_rom[61][51] = 8'd202;
	sample_rom[61][52] = 8'd199;
	sample_rom[61][53] = 8'd197;
	sample_rom[61][54] = 8'd192;
	sample_rom[61][55] = 8'd187;
	sample_rom[61][56] = 8'd182;
	sample_rom[61][57] = 8'd176;
	sample_rom[61][58] = 8'd169;
	sample_rom[61][59] = 8'd164;
	sample_rom[61][60] = 8'd157;
	sample_rom[61][61] = 8'd149;
	sample_rom[61][62] = 8'd141;
	sample_rom[61][63] = 8'd133;
	sample_rom[62][0] = 8'd129;
	sample_rom[62][1] = 8'd142;
	sample_rom[62][2] = 8'd153;
	sample_rom[62][3] = 8'd162;
	sample_rom[62][4] = 8'd171;
	sample_rom[62][5] = 8'd181;
	sample_rom[62][6] = 8'd188;
	sample_rom[62][7] = 8'd196;
	sample_rom[62][8] = 8'd201;
	sample_rom[62][9] = 8'd207;
	sample_rom[62][10] = 8'd212;
	sample_rom[62][11] = 8'd214;
	sample_rom[62][12] = 8'd216;
	sample_rom[62][13] = 8'd218;
	sample_rom[62][14] = 8'd220;
	sample_rom[62][15] = 8'd220;
	sample_rom[62][16] = 8'd219;
	sample_rom[62][17] = 8'd217;
	sample_rom[62][18] = 8'd214;
	sample_rom[62][19] = 8'd210;
	sample_rom[62][20] = 8'd207;
	sample_rom[62][21] = 8'd202;
	sample_rom[62][22] = 8'd195;
	sample_rom[62][23] = 8'd192;
	sample_rom[62][24] = 8'd186;
	sample_rom[62][25] = 8'd180;
	sample_rom[62][26] = 8'd171;
	sample_rom[62][27] = 8'd165;
	sample_rom[62][28] = 8'd160;
	sample_rom[62][29] = 8'd155;
	sample_rom[62][30] = 8'd149;
	sample_rom[62][31] = 8'd141;
	sample_rom[62][32] = 8'd136;
	sample_rom[62][33] = 8'd129;
	sample_rom[62][34] = 8'd123;
	sample_rom[62][35] = 8'd122;
	sample_rom[62][36] = 8'd119;
	sample_rom[62][37] = 8'd113;
	sample_rom[62][38] = 8'd110;
	sample_rom[62][39] = 8'd107;
	sample_rom[62][40] = 8'd106;
	sample_rom[62][41] = 8'd103;
	sample_rom[62][42] = 8'd104;
	sample_rom[62][43] = 8'd102;
	sample_rom[62][44] = 8'd103;
	sample_rom[62][45] = 8'd101;
	sample_rom[62][46] = 8'd101;
	sample_rom[62][47] = 8'd101;
	sample_rom[62][48] = 8'd101;
	sample_rom[62][49] = 8'd104;
	sample_rom[62][50] = 8'd105;
	sample_rom[62][51] = 8'd105;
	sample_rom[62][52] = 8'd108;
	sample_rom[62][53] = 8'd109;
	sample_rom[62][54] = 8'd114;
	sample_rom[62][55] = 8'd113;
	sample_rom[62][56] = 8'd115;
	sample_rom[62][57] = 8'd119;
	sample_rom[62][58] = 8'd121;
	sample_rom[62][59] = 8'd123;
	sample_rom[62][60] = 8'd124;
	sample_rom[62][61] = 8'd127;
	sample_rom[62][62] = 8'd125;
	sample_rom[62][63] = 8'd127;
	sample_rom[63][0] = 8'd129;
	sample_rom[63][1] = 8'd142;
	sample_rom[63][2] = 8'd152;
	sample_rom[63][3] = 8'd160;
	sample_rom[63][4] = 8'd168;
	sample_rom[63][5] = 8'd178;
	sample_rom[63][6] = 8'd185;
	sample_rom[63][7] = 8'd193;
	sample_rom[63][8] = 8'd199;
	sample_rom[63][9] = 8'd205;
	sample_rom[63][10] = 8'd210;
	sample_rom[63][11] = 8'd214;
	sample_rom[63][12] = 8'd216;
	sample_rom[63][13] = 8'd218;
	sample_rom[63][14] = 8'd221;
	sample_rom[63][15] = 8'd221;
	sample_rom[63][16] = 8'd221;
	sample_rom[63][17] = 8'd218;
	sample_rom[63][18] = 8'd215;
	sample_rom[63][19] = 8'd212;
	sample_rom[63][20] = 8'd208;
	sample_rom[63][21] = 8'd203;
	sample_rom[63][22] = 8'd196;
	sample_rom[63][23] = 8'd193;
	sample_rom[63][24] = 8'd186;
	sample_rom[63][25] = 8'd180;
	sample_rom[63][26] = 8'd172;
	sample_rom[63][27] = 8'd166;
	sample_rom[63][28] = 8'd160;
	sample_rom[63][29] = 8'd154;
	sample_rom[63][30] = 8'd149;
	sample_rom[63][31] = 8'd141;
	sample_rom[63][32] = 8'd136;
	sample_rom[63][33] = 8'd129;
	sample_rom[63][34] = 8'd123;
	sample_rom[63][35] = 8'd120;
	sample_rom[63][36] = 8'd117;
	sample_rom[63][37] = 8'd112;
	sample_rom[63][38] = 8'd109;
	sample_rom[63][39] = 8'd105;
	sample_rom[63][40] = 8'd104;
	sample_rom[63][41] = 8'd102;
	sample_rom[63][42] = 8'd103;
	sample_rom[63][43] = 8'd101;
	sample_rom[63][44] = 8'd102;
	sample_rom[63][45] = 8'd101;
	sample_rom[63][46] = 8'd102;
	sample_rom[63][47] = 8'd102;
	sample_rom[63][48] = 8'd103;
	sample_rom[63][49] = 8'd105;
	sample_rom[63][50] = 8'd106;
	sample_rom[63][51] = 8'd107;
	sample_rom[63][52] = 8'd110;
	sample_rom[63][53] = 8'd111;
	sample_rom[63][54] = 8'd114;
	sample_rom[63][55] = 8'd113;
	sample_rom[63][56] = 8'd115;
	sample_rom[63][57] = 8'd118;
	sample_rom[63][58] = 8'd120;
	sample_rom[63][59] = 8'd122;
	sample_rom[63][60] = 8'd123;
	sample_rom[63][61] = 8'd125;
	sample_rom[63][62] = 8'd124;
	sample_rom[63][63] = 8'd127;
	sample_rom[64][0] = 8'd130;
	sample_rom[64][1] = 8'd148;
	sample_rom[64][2] = 8'd164;
	sample_rom[64][3] = 8'd178;
	sample_rom[64][4] = 8'd192;
	sample_rom[64][5] = 8'd205;
	sample_rom[64][6] = 8'd215;
	sample_rom[64][7] = 8'd223;
	sample_rom[64][8] = 8'd47;
	sample_rom[64][9] = 8'd255;
	sample_rom[64][10] = 8'd236;
	sample_rom[64][11] = 8'd236;
	sample_rom[64][12] = 8'd237;
	sample_rom[64][13] = 8'd235;
	sample_rom[64][14] = 8'd231;
	sample_rom[64][15] = 8'd228;
	sample_rom[64][16] = 8'd223;
	sample_rom[64][17] = 8'd217;
	sample_rom[64][18] = 8'd210;
	sample_rom[64][19] = 8'd205;
	sample_rom[64][20] = 8'd199;
	sample_rom[64][21] = 8'd195;
	sample_rom[64][22] = 8'd189;
	sample_rom[64][23] = 8'd186;
	sample_rom[64][24] = 8'd182;
	sample_rom[64][25] = 8'd180;
	sample_rom[64][26] = 8'd178;
	sample_rom[64][27] = 8'd177;
	sample_rom[64][28] = 8'd176;
	sample_rom[64][29] = 8'd174;
	sample_rom[64][30] = 8'd175;
	sample_rom[64][31] = 8'd174;
	sample_rom[64][32] = 8'd172;
	sample_rom[64][33] = 8'd171;
	sample_rom[64][34] = 8'd168;
	sample_rom[64][35] = 8'd167;
	sample_rom[64][36] = 8'd162;
	sample_rom[64][37] = 8'd160;
	sample_rom[64][38] = 8'd156;
	sample_rom[64][39] = 8'd149;
	sample_rom[64][40] = 8'd146;
	sample_rom[64][41] = 8'd139;
	sample_rom[64][42] = 8'd135;
	sample_rom[64][43] = 8'd128;
	sample_rom[64][44] = 8'd122;
	sample_rom[64][45] = 8'd116;
	sample_rom[64][46] = 8'd111;
	sample_rom[64][47] = 8'd105;
	sample_rom[64][48] = 8'd101;
	sample_rom[64][49] = 8'd98;
	sample_rom[64][50] = 8'd96;
	sample_rom[64][51] = 8'd94;
	sample_rom[64][52] = 8'd93;
	sample_rom[64][53] = 8'd93;
	sample_rom[64][54] = 8'd94;
	sample_rom[64][55] = 8'd95;
	sample_rom[64][56] = 8'd96;
	sample_rom[64][57] = 8'd99;
	sample_rom[64][58] = 8'd102;
	sample_rom[64][59] = 8'd106;
	sample_rom[64][60] = 8'd108;
	sample_rom[64][61] = 8'd114;
	sample_rom[64][62] = 8'd118;
	sample_rom[64][63] = 8'd124;
	sample_rom[65][0] = 8'd130;
	sample_rom[65][1] = 8'd140;
	sample_rom[65][2] = 8'd151;
	sample_rom[65][3] = 8'd160;
	sample_rom[65][4] = 8'd169;
	sample_rom[65][5] = 8'd176;
	sample_rom[65][6] = 8'd185;
	sample_rom[65][7] = 8'd193;
	sample_rom[65][8] = 8'd199;
	sample_rom[65][9] = 8'd207;
	sample_rom[65][10] = 8'd212;
	sample_rom[65][11] = 8'd218;
	sample_rom[65][12] = 8'd223;
	sample_rom[65][13] = 8'd225;
	sample_rom[65][14] = 8'd229;
	sample_rom[65][15] = 8'd232;
	sample_rom[65][16] = 8'd234;
	sample_rom[65][17] = 8'd235;
	sample_rom[65][18] = 8'd236;
	sample_rom[65][19] = 8'd236;
	sample_rom[65][20] = 8'd233;
	sample_rom[65][21] = 8'd233;
	sample_rom[65][22] = 8'd230;
	sample_rom[65][23] = 8'd228;
	sample_rom[65][24] = 8'd225;
	sample_rom[65][25] = 8'd223;
	sample_rom[65][26] = 8'd218;
	sample_rom[65][27] = 8'd214;
	sample_rom[65][28] = 8'd210;
	sample_rom[65][29] = 8'd206;
	sample_rom[65][30] = 8'd201;
	sample_rom[65][31] = 8'd195;
	sample_rom[65][32] = 8'd191;
	sample_rom[65][33] = 8'd186;
	sample_rom[65][34] = 8'd181;
	sample_rom[65][35] = 8'd177;
	sample_rom[65][36] = 8'd172;
	sample_rom[65][37] = 8'd167;
	sample_rom[65][38] = 8'd164;
	sample_rom[65][39] = 8'd160;
	sample_rom[65][40] = 8'd156;
	sample_rom[65][41] = 8'd152;
	sample_rom[65][42] = 8'd150;
	sample_rom[65][43] = 8'd146;
	sample_rom[65][44] = 8'd144;
	sample_rom[65][45] = 8'd142;
	sample_rom[65][46] = 8'd139;
	sample_rom[65][47] = 8'd137;
	sample_rom[65][48] = 8'd136;
	sample_rom[65][49] = 8'd133;
	sample_rom[65][50] = 8'd132;
	sample_rom[65][51] = 8'd131;
	sample_rom[65][52] = 8'd130;
	sample_rom[65][53] = 8'd129;
	sample_rom[65][54] = 8'd129;
	sample_rom[65][55] = 8'd128;
	sample_rom[65][56] = 8'd128;
	sample_rom[65][57] = 8'd127;
	sample_rom[65][58] = 8'd127;
	sample_rom[65][59] = 8'd128;
	sample_rom[65][60] = 8'd127;
	sample_rom[65][61] = 8'd127;
	sample_rom[65][62] = 8'd126;
	sample_rom[65][63] = 8'd127;
	sample_rom[66][0] = 8'd132;
	sample_rom[66][1] = 8'd170;
	sample_rom[66][2] = 8'd202;
	sample_rom[66][3] = 8'd230;
	sample_rom[66][4] = 8'd245;
	sample_rom[66][5] = 8'd253;
	sample_rom[66][6] = 8'd253;
	sample_rom[66][7] = 8'd246;
	sample_rom[66][8] = 8'd236;
	sample_rom[66][9] = 8'd227;
	sample_rom[66][10] = 8'd216;
	sample_rom[66][11] = 8'd206;
	sample_rom[66][12] = 8'd195;
	sample_rom[66][13] = 8'd183;
	sample_rom[66][14] = 8'd173;
	sample_rom[66][15] = 8'd158;
	sample_rom[66][16] = 8'd144;
	sample_rom[66][17] = 8'd131;
	sample_rom[66][18] = 8'd123;
	sample_rom[66][19] = 8'd113;
	sample_rom[66][20] = 8'd108;
	sample_rom[66][21] = 8'd108;
	sample_rom[66][22] = 8'd110;
	sample_rom[66][23] = 8'd119;
	sample_rom[66][24] = 8'd124;
	sample_rom[66][25] = 8'd127;
	sample_rom[66][26] = 8'd131;
	sample_rom[66][27] = 8'd139;
	sample_rom[66][28] = 8'd145;
	sample_rom[66][29] = 8'd155;
	sample_rom[66][30] = 8'd166;
	sample_rom[66][31] = 8'd177;
	sample_rom[66][32] = 8'd188;
	sample_rom[66][33] = 8'd201;
	sample_rom[66][34] = 8'd207;
	sample_rom[66][35] = 8'd211;
	sample_rom[66][36] = 8'd210;
	sample_rom[66][37] = 8'd200;
	sample_rom[66][38] = 8'd190;
	sample_rom[66][39] = 8'd176;
	sample_rom[66][40] = 8'd164;
	sample_rom[66][41] = 8'd153;
	sample_rom[66][42] = 8'd143;
	sample_rom[66][43] = 8'd135;
	sample_rom[66][44] = 8'd129;
	sample_rom[66][45] = 8'd127;
	sample_rom[66][46] = 8'd121;
	sample_rom[66][47] = 8'd116;
	sample_rom[66][48] = 8'd110;
	sample_rom[66][49] = 8'd107;
	sample_rom[66][50] = 8'd103;
	sample_rom[66][51] = 8'd100;
	sample_rom[66][52] = 8'd103;
	sample_rom[66][53] = 8'd106;
	sample_rom[66][54] = 8'd112;
	sample_rom[66][55] = 8'd118;
	sample_rom[66][56] = 8'd122;
	sample_rom[66][57] = 8'd127;
	sample_rom[66][58] = 8'd130;
	sample_rom[66][59] = 8'd133;
	sample_rom[66][60] = 8'd132;
	sample_rom[66][61] = 8'd131;
	sample_rom[66][62] = 8'd130;
	sample_rom[66][63] = 8'd128;
	sample_rom[67][0] = 8'd132;
	sample_rom[67][1] = 8'd183;
	sample_rom[67][2] = 8'd223;
	sample_rom[67][3] = 8'd246;
	sample_rom[67][4] = 8'd245;
	sample_rom[67][5] = 8'd223;
	sample_rom[67][6] = 8'd188;
	sample_rom[67][7] = 8'd143;
	sample_rom[67][8] = 8'd100;
	sample_rom[67][9] = 8'd70;
	sample_rom[67][10] = 8'd52;
	sample_rom[67][11] = 8'd56;
	sample_rom[67][12] = 8'd76;
	sample_rom[67][13] = 8'd107;
	sample_rom[67][14] = 8'd148;
	sample_rom[67][15] = 8'd185;
	sample_rom[67][16] = 8'd215;
	sample_rom[67][17] = 8'd233;
	sample_rom[67][18] = 8'd236;
	sample_rom[67][19] = 8'd223;
	sample_rom[67][20] = 8'd203;
	sample_rom[67][21] = 8'd174;
	sample_rom[67][22] = 8'd142;
	sample_rom[67][23] = 8'd116;
	sample_rom[67][24] = 8'd97;
	sample_rom[67][25] = 8'd91;
	sample_rom[67][26] = 8'd97;
	sample_rom[67][27] = 8'd115;
	sample_rom[67][28] = 8'd140;
	sample_rom[67][29] = 8'd166;
	sample_rom[67][30] = 8'd192;
	sample_rom[67][31] = 8'd206;
	sample_rom[67][32] = 8'd210;
	sample_rom[67][33] = 8'd201;
	sample_rom[67][34] = 8'd182;
	sample_rom[67][35] = 8'd161;
	sample_rom[67][36] = 8'd141;
	sample_rom[67][37] = 8'd121;
	sample_rom[67][38] = 8'd111;
	sample_rom[67][39] = 8'd108;
	sample_rom[67][40] = 8'd112;
	sample_rom[67][41] = 8'd121;
	sample_rom[67][42] = 8'd137;
	sample_rom[67][43] = 8'd147;
	sample_rom[67][44] = 8'd156;
	sample_rom[67][45] = 8'd161;
	sample_rom[67][46] = 8'd163;
	sample_rom[67][47] = 8'd159;
	sample_rom[67][48] = 8'd156;
	sample_rom[67][49] = 8'd147;
	sample_rom[67][50] = 8'd141;
	sample_rom[67][51] = 8'd131;
	sample_rom[67][52] = 8'd124;
	sample_rom[67][53] = 8'd117;
	sample_rom[67][54] = 8'd113;
	sample_rom[67][55] = 8'd111;
	sample_rom[67][56] = 8'd117;
	sample_rom[67][57] = 8'd125;
	sample_rom[67][58] = 8'd134;
	sample_rom[67][59] = 8'd143;
	sample_rom[67][60] = 8'd149;
	sample_rom[67][61] = 8'd150;
	sample_rom[67][62] = 8'd147;
	sample_rom[67][63] = 8'd138;
	sample_rom[68][0] = 8'd132;
	sample_rom[68][1] = 8'd199;
	sample_rom[68][2] = 8'd228;
	sample_rom[68][3] = 8'd211;
	sample_rom[68][4] = 8'd151;
	sample_rom[68][5] = 8'd86;
	sample_rom[68][6] = 8'd52;
	sample_rom[68][7] = 8'd66;
	sample_rom[68][8] = 8'd118;
	sample_rom[68][9] = 8'd184;
	sample_rom[68][10] = 8'd226;
	sample_rom[68][11] = 8'd226;
	sample_rom[68][12] = 8'd186;
	sample_rom[68][13] = 8'd130;
	sample_rom[68][14] = 8'd91;
	sample_rom[68][15] = 8'd86;
	sample_rom[68][16] = 8'd116;
	sample_rom[68][17] = 8'd164;
	sample_rom[68][18] = 8'd205;
	sample_rom[68][19] = 8'd214;
	sample_rom[68][20] = 8'd195;
	sample_rom[68][21] = 8'd160;
	sample_rom[68][22] = 8'd126;
	sample_rom[68][23] = 8'd114;
	sample_rom[68][24] = 8'd125;
	sample_rom[68][25] = 8'd153;
	sample_rom[68][26] = 8'd177;
	sample_rom[68][27] = 8'd188;
	sample_rom[68][28] = 8'd180;
	sample_rom[68][29] = 8'd162;
	sample_rom[68][30] = 8'd146;
	sample_rom[68][31] = 8'd137;
	sample_rom[68][32] = 8'd138;
	sample_rom[68][33] = 8'd147;
	sample_rom[68][34] = 8'd157;
	sample_rom[68][35] = 8'd160;
	sample_rom[68][36] = 8'd159;
	sample_rom[68][37] = 8'd151;
	sample_rom[68][38] = 8'd145;
	sample_rom[68][39] = 8'd142;
	sample_rom[68][40] = 8'd145;
	sample_rom[68][41] = 8'd145;
	sample_rom[68][42] = 8'd146;
	sample_rom[68][43] = 8'd142;
	sample_rom[68][44] = 8'd138;
	sample_rom[68][45] = 8'd138;
	sample_rom[68][46] = 8'd137;
	sample_rom[68][47] = 8'd139;
	sample_rom[68][48] = 8'd142;
	sample_rom[68][49] = 8'd141;
	sample_rom[68][50] = 8'd140;
	sample_rom[68][51] = 8'd135;
	sample_rom[68][52] = 8'd130;
	sample_rom[68][53] = 8'd127;
	sample_rom[68][54] = 8'd128;
	sample_rom[68][55] = 8'd131;
	sample_rom[68][56] = 8'd136;
	sample_rom[68][57] = 8'd137;
	sample_rom[68][58] = 8'd134;
	sample_rom[68][59] = 8'd132;
	sample_rom[68][60] = 8'd128;
	sample_rom[68][61] = 8'd124;
	sample_rom[68][62] = 8'd123;
	sample_rom[68][63] = 8'd125;
	sample_rom[69][0] = 8'd130;
	sample_rom[69][1] = 8'd139;
	sample_rom[69][2] = 8'd148;
	sample_rom[69][3] = 8'd154;
	sample_rom[69][4] = 8'd161;
	sample_rom[69][5] = 8'd169;
	sample_rom[69][6] = 8'd175;
	sample_rom[69][7] = 8'd182;
	sample_rom[69][8] = 8'd189;
	sample_rom[69][9] = 8'd194;
	sample_rom[69][10] = 8'd199;
	sample_rom[69][11] = 8'd204;
	sample_rom[69][12] = 8'd208;
	sample_rom[69][13] = 8'd211;
	sample_rom[69][14] = 8'd215;
	sample_rom[69][15] = 8'd218;
	sample_rom[69][16] = 8'd219;
	sample_rom[69][17] = 8'd220;
	sample_rom[69][18] = 8'd220;
	sample_rom[69][19] = 8'd220;
	sample_rom[69][20] = 8'd218;
	sample_rom[69][21] = 8'd217;
	sample_rom[69][22] = 8'd214;
	sample_rom[69][23] = 8'd213;
	sample_rom[69][24] = 8'd210;
	sample_rom[69][25] = 8'd206;
	sample_rom[69][26] = 8'd201;
	sample_rom[69][27] = 8'd197;
	sample_rom[69][28] = 8'd191;
	sample_rom[69][29] = 8'd187;
	sample_rom[69][30] = 8'd182;
	sample_rom[69][31] = 8'd175;
	sample_rom[69][32] = 8'd170;
	sample_rom[69][33] = 8'd163;
	sample_rom[69][34] = 8'd158;
	sample_rom[69][35] = 8'd153;
	sample_rom[69][36] = 8'd147;
	sample_rom[69][37] = 8'd140;
	sample_rom[69][38] = 8'd136;
	sample_rom[69][39] = 8'd130;
	sample_rom[69][40] = 8'd124;
	sample_rom[69][41] = 8'd121;
	sample_rom[69][42] = 8'd116;
	sample_rom[69][43] = 8'd112;
	sample_rom[69][44] = 8'd109;
	sample_rom[69][45] = 8'd106;
	sample_rom[69][46] = 8'd103;
	sample_rom[69][47] = 8'd100;
	sample_rom[69][48] = 8'd99;
	sample_rom[69][49] = 8'd98;
	sample_rom[69][50] = 8'd97;
	sample_rom[69][51] = 8'd97;
	sample_rom[69][52] = 8'd98;
	sample_rom[69][53] = 8'd98;
	sample_rom[69][54] = 8'd100;
	sample_rom[69][55] = 8'd101;
	sample_rom[69][56] = 8'd102;
	sample_rom[69][57] = 8'd105;
	sample_rom[69][58] = 8'd108;
	sample_rom[69][59] = 8'd111;
	sample_rom[69][60] = 8'd115;
	sample_rom[69][61] = 8'd119;
	sample_rom[69][62] = 8'd120;
	sample_rom[69][63] = 8'd125;
	sample_rom[70][0] = 8'd130;
	sample_rom[70][1] = 8'd142;
	sample_rom[70][2] = 8'd154;
	sample_rom[70][3] = 8'd163;
	sample_rom[70][4] = 8'd173;
	sample_rom[70][5] = 8'd182;
	sample_rom[70][6] = 8'd190;
	sample_rom[70][7] = 8'd198;
	sample_rom[70][8] = 8'd203;
	sample_rom[70][9] = 8'd209;
	sample_rom[70][10] = 8'd214;
	sample_rom[70][11] = 8'd216;
	sample_rom[70][12] = 8'd216;
	sample_rom[70][13] = 8'd216;
	sample_rom[70][14] = 8'd215;
	sample_rom[70][15] = 8'd212;
	sample_rom[70][16] = 8'd209;
	sample_rom[70][17] = 8'd204;
	sample_rom[70][18] = 8'd198;
	sample_rom[70][19] = 8'd192;
	sample_rom[70][20] = 8'd185;
	sample_rom[70][21] = 8'd178;
	sample_rom[70][22] = 8'd171;
	sample_rom[70][23] = 8'd165;
	sample_rom[70][24] = 8'd158;
	sample_rom[70][25] = 8'd152;
	sample_rom[70][26] = 8'd145;
	sample_rom[70][27] = 8'd140;
	sample_rom[70][28] = 8'd137;
	sample_rom[70][29] = 8'd133;
	sample_rom[70][30] = 8'd131;
	sample_rom[70][31] = 8'd129;
	sample_rom[70][32] = 8'd128;
	sample_rom[70][33] = 8'd129;
	sample_rom[70][34] = 8'd130;
	sample_rom[70][35] = 8'd134;
	sample_rom[70][36] = 8'd137;
	sample_rom[70][37] = 8'd141;
	sample_rom[70][38] = 8'd147;
	sample_rom[70][39] = 8'd152;
	sample_rom[70][40] = 8'd160;
	sample_rom[70][41] = 8'd165;
	sample_rom[70][42] = 8'd173;
	sample_rom[70][43] = 8'd179;
	sample_rom[70][44] = 8'd187;
	sample_rom[70][45] = 8'd193;
	sample_rom[70][46] = 8'd200;
	sample_rom[70][47] = 8'd205;
	sample_rom[70][48] = 8'd209;
	sample_rom[70][49] = 8'd212;
	sample_rom[70][50] = 8'd214;
	sample_rom[70][51] = 8'd215;
	sample_rom[70][52] = 8'd215;
	sample_rom[70][53] = 8'd214;
	sample_rom[70][54] = 8'd210;
	sample_rom[70][55] = 8'd205;
	sample_rom[70][56] = 8'd201;
	sample_rom[70][57] = 8'd193;
	sample_rom[70][58] = 8'd186;
	sample_rom[70][59] = 8'd178;
	sample_rom[70][60] = 8'd168;
	sample_rom[70][61] = 8'd159;
	sample_rom[70][62] = 8'd147;
	sample_rom[70][63] = 8'd137;
	sample_rom[71][0] = 8'd130;
	sample_rom[71][1] = 8'd145;
	sample_rom[71][2] = 8'd159;
	sample_rom[71][3] = 8'd170;
	sample_rom[71][4] = 8'd182;
	sample_rom[71][5] = 8'd190;
	sample_rom[71][6] = 8'd198;
	sample_rom[71][7] = 8'd205;
	sample_rom[71][8] = 8'd208;
	sample_rom[71][9] = 8'd209;
	sample_rom[71][10] = 8'd209;
	sample_rom[71][11] = 8'd205;
	sample_rom[71][12] = 8'd200;
	sample_rom[71][13] = 8'd194;
	sample_rom[71][14] = 8'd186;
	sample_rom[71][15] = 8'd177;
	sample_rom[71][16] = 8'd168;
	sample_rom[71][17] = 8'd159;
	sample_rom[71][18] = 8'd150;
	sample_rom[71][19] = 8'd142;
	sample_rom[71][20] = 8'd134;
	sample_rom[71][21] = 8'd130;
	sample_rom[71][22] = 8'd126;
	sample_rom[71][23] = 8'd124;
	sample_rom[71][24] = 8'd123;
	sample_rom[71][25] = 8'd127;
	sample_rom[71][26] = 8'd131;
	sample_rom[71][27] = 8'd137;
	sample_rom[71][28] = 8'd145;
	sample_rom[71][29] = 8'd154;
	sample_rom[71][30] = 8'd164;
	sample_rom[71][31] = 8'd175;
	sample_rom[71][32] = 8'd186;
	sample_rom[71][33] = 8'd198;
	sample_rom[71][34] = 8'd207;
	sample_rom[71][35] = 8'd217;
	sample_rom[71][36] = 8'd224;
	sample_rom[71][37] = 8'd229;
	sample_rom[71][38] = 8'd234;
	sample_rom[71][39] = 8'd236;
	sample_rom[71][40] = 8'd237;
	sample_rom[71][41] = 8'd233;
	sample_rom[71][42] = 8'd229;
	sample_rom[71][43] = 8'd222;
	sample_rom[71][44] = 8'd214;
	sample_rom[71][45] = 8'd203;
	sample_rom[71][46] = 8'd192;
	sample_rom[71][47] = 8'd179;
	sample_rom[71][48] = 8'd166;
	sample_rom[71][49] = 8'd153;
	sample_rom[71][50] = 8'd141;
	sample_rom[71][51] = 8'd128;
	sample_rom[71][52] = 8'd117;
	sample_rom[71][53] = 8'd109;
	sample_rom[71][54] = 8'd101;
	sample_rom[71][55] = 8'd95;
	sample_rom[71][56] = 8'd92;
	sample_rom[71][57] = 8'd91;
	sample_rom[71][58] = 8'd92;
	sample_rom[71][59] = 8'd95;
	sample_rom[71][60] = 8'd98;
	sample_rom[71][61] = 8'd105;
	sample_rom[71][62] = 8'd111;
	sample_rom[71][63] = 8'd119;
	sample_rom[72][0] = 8'd130;
	sample_rom[72][1] = 8'd147;
	sample_rom[72][2] = 8'd164;
	sample_rom[72][3] = 8'd177;
	sample_rom[72][4] = 8'd188;
	sample_rom[72][5] = 8'd197;
	sample_rom[72][6] = 8'd203;
	sample_rom[72][7] = 8'd205;
	sample_rom[72][8] = 8'd203;
	sample_rom[72][9] = 8'd198;
	sample_rom[72][10] = 8'd192;
	sample_rom[72][11] = 8'd181;
	sample_rom[72][12] = 8'd170;
	sample_rom[72][13] = 8'd160;
	sample_rom[72][14] = 8'd148;
	sample_rom[72][15] = 8'd137;
	sample_rom[72][16] = 8'd128;
	sample_rom[72][17] = 8'd122;
	sample_rom[72][18] = 8'd118;
	sample_rom[72][19] = 8'd117;
	sample_rom[72][20] = 8'd120;
	sample_rom[72][21] = 8'd127;
	sample_rom[72][22] = 8'd135;
	sample_rom[72][23] = 8'd148;
	sample_rom[72][24] = 8'd160;
	sample_rom[72][25] = 8'd175;
	sample_rom[72][26] = 8'd190;
	sample_rom[72][27] = 8'd204;
	sample_rom[72][28] = 8'd217;
	sample_rom[72][29] = 8'd227;
	sample_rom[72][30] = 8'd235;
	sample_rom[72][31] = 8'd240;
	sample_rom[72][32] = 8'd242;
	sample_rom[72][33] = 8'd239;
	sample_rom[72][34] = 8'd233;
	sample_rom[72][35] = 8'd225;
	sample_rom[72][36] = 8'd214;
	sample_rom[72][37] = 8'd200;
	sample_rom[72][38] = 8'd186;
	sample_rom[72][39] = 8'd170;
	sample_rom[72][40] = 8'd158;
	sample_rom[72][41] = 8'd143;
	sample_rom[72][42] = 8'd133;
	sample_rom[72][43] = 8'd124;
	sample_rom[72][44] = 8'd118;
	sample_rom[72][45] = 8'd115;
	sample_rom[72][46] = 8'd117;
	sample_rom[72][47] = 8'd122;
	sample_rom[72][48] = 8'd128;
	sample_rom[72][49] = 8'd137;
	sample_rom[72][50] = 8'd149;
	sample_rom[72][51] = 8'd160;
	sample_rom[72][52] = 8'd171;
	sample_rom[72][53] = 8'd182;
	sample_rom[72][54] = 8'd191;
	sample_rom[72][55] = 8'd197;
	sample_rom[72][56] = 8'd201;
	sample_rom[72][57] = 8'd202;
	sample_rom[72][58] = 8'd199;
	sample_rom[72][59] = 8'd193;
	sample_rom[72][60] = 8'd184;
	sample_rom[72][61] = 8'd173;
	sample_rom[72][62] = 8'd158;
	sample_rom[72][63] = 8'd142;
	sample_rom[73][0] = 8'd130;
	sample_rom[73][1] = 8'd150;
	sample_rom[73][2] = 8'd168;
	sample_rom[73][3] = 8'd182;
	sample_rom[73][4] = 8'd193;
	sample_rom[73][5] = 8'd200;
	sample_rom[73][6] = 8'd201;
	sample_rom[73][7] = 8'd198;
	sample_rom[73][8] = 8'd190;
	sample_rom[73][9] = 8'd179;
	sample_rom[73][10] = 8'd166;
	sample_rom[73][11] = 8'd152;
	sample_rom[73][12] = 8'd138;
	sample_rom[73][13] = 8'd126;
	sample_rom[73][14] = 8'd118;
	sample_rom[73][15] = 8'd113;
	sample_rom[73][16] = 8'd112;
	sample_rom[73][17] = 8'd117;
	sample_rom[73][18] = 8'd126;
	sample_rom[73][19] = 8'd139;
	sample_rom[73][20] = 8'd155;
	sample_rom[73][21] = 8'd173;
	sample_rom[73][22] = 8'd191;
	sample_rom[73][23] = 8'd209;
	sample_rom[73][24] = 8'd222;
	sample_rom[73][25] = 8'd232;
	sample_rom[73][26] = 8'd238;
	sample_rom[73][27] = 8'd239;
	sample_rom[73][28] = 8'd236;
	sample_rom[73][29] = 8'd227;
	sample_rom[73][30] = 8'd216;
	sample_rom[73][31] = 8'd200;
	sample_rom[73][32] = 8'd184;
	sample_rom[73][33] = 8'd167;
	sample_rom[73][34] = 8'd152;
	sample_rom[73][35] = 8'd140;
	sample_rom[73][36] = 8'd131;
	sample_rom[73][37] = 8'd125;
	sample_rom[73][38] = 8'd127;
	sample_rom[73][39] = 8'd131;
	sample_rom[73][40] = 8'd141;
	sample_rom[73][41] = 8'd153;
	sample_rom[73][42] = 8'd167;
	sample_rom[73][43] = 8'd183;
	sample_rom[73][44] = 8'd197;
	sample_rom[73][45] = 8'd210;
	sample_rom[73][46] = 8'd219;
	sample_rom[73][47] = 8'd223;
	sample_rom[73][48] = 8'd224;
	sample_rom[73][49] = 8'd220;
	sample_rom[73][50] = 8'd210;
	sample_rom[73][51] = 8'd196;
	sample_rom[73][52] = 8'd179;
	sample_rom[73][53] = 8'd160;
	sample_rom[73][54] = 8'd141;
	sample_rom[73][55] = 8'd122;
	sample_rom[73][56] = 8'd107;
	sample_rom[73][57] = 8'd96;
	sample_rom[73][58] = 8'd87;
	sample_rom[73][59] = 8'd85;
	sample_rom[73][60] = 8'd87;
	sample_rom[73][61] = 8'd93;
	sample_rom[73][62] = 8'd101;
	sample_rom[73][63] = 8'd114;
	sample_rom[74][0] = 8'd130;
	sample_rom[74][1] = 8'd157;
	sample_rom[74][2] = 8'd181;
	sample_rom[74][3] = 8'd197;
	sample_rom[74][4] = 8'd209;
	sample_rom[74][5] = 8'd209;
	sample_rom[74][6] = 8'd203;
	sample_rom[74][7] = 8'd190;
	sample_rom[74][8] = 8'd173;
	sample_rom[74][9] = 8'd153;
	sample_rom[74][10] = 8'd134;
	sample_rom[74][11] = 8'd117;
	sample_rom[74][12] = 8'd104;
	sample_rom[74][13] = 8'd100;
	sample_rom[74][14] = 8'd103;
	sample_rom[74][15] = 8'd113;
	sample_rom[74][16] = 8'd128;
	sample_rom[74][17] = 8'd149;
	sample_rom[74][18] = 8'd170;
	sample_rom[74][19] = 8'd192;
	sample_rom[74][20] = 8'd212;
	sample_rom[74][21] = 8'd227;
	sample_rom[74][22] = 8'd235;
	sample_rom[74][23] = 8'd239;
	sample_rom[74][24] = 8'd234;
	sample_rom[74][25] = 8'd224;
	sample_rom[74][26] = 8'd208;
	sample_rom[74][27] = 8'd191;
	sample_rom[74][28] = 8'd171;
	sample_rom[74][29] = 8'd154;
	sample_rom[74][30] = 8'd141;
	sample_rom[74][31] = 8'd131;
	sample_rom[74][32] = 8'd128;
	sample_rom[74][33] = 8'd133;
	sample_rom[74][34] = 8'd141;
	sample_rom[74][35] = 8'd156;
	sample_rom[74][36] = 8'd173;
	sample_rom[74][37] = 8'd192;
	sample_rom[74][38] = 8'd211;
	sample_rom[74][39] = 8'd223;
	sample_rom[74][40] = 8'd230;
	sample_rom[74][41] = 8'd233;
	sample_rom[74][42] = 8'd228;
	sample_rom[74][43] = 8'd217;
	sample_rom[74][44] = 8'd202;
	sample_rom[74][45] = 8'd183;
	sample_rom[74][46] = 8'd162;
	sample_rom[74][47] = 8'd144;
	sample_rom[74][48] = 8'd128;
	sample_rom[74][49] = 8'd118;
	sample_rom[74][50] = 8'd112;
	sample_rom[74][51] = 8'd113;
	sample_rom[74][52] = 8'd120;
	sample_rom[74][53] = 8'd131;
	sample_rom[74][54] = 8'd144;
	sample_rom[74][55] = 8'd157;
	sample_rom[74][56] = 8'd169;
	sample_rom[74][57] = 8'd181;
	sample_rom[74][58] = 8'd185;
	sample_rom[74][59] = 8'd187;
	sample_rom[74][60] = 8'd182;
	sample_rom[74][61] = 8'd173;
	sample_rom[74][62] = 8'd160;
	sample_rom[74][63] = 8'd143;
	sample_rom[75][0] = 8'd130;
	sample_rom[75][1] = 8'd160;
	sample_rom[75][2] = 8'd187;
	sample_rom[75][3] = 8'd201;
	sample_rom[75][4] = 8'd210;
	sample_rom[75][5] = 8'd205;
	sample_rom[75][6] = 8'd191;
	sample_rom[75][7] = 8'd171;
	sample_rom[75][8] = 8'd147;
	sample_rom[75][9] = 8'd125;
	sample_rom[75][10] = 8'd107;
	sample_rom[75][11] = 8'd97;
	sample_rom[75][12] = 8'd96;
	sample_rom[75][13] = 8'd106;
	sample_rom[75][14] = 8'd124;
	sample_rom[75][15] = 8'd148;
	sample_rom[75][16] = 8'd172;
	sample_rom[75][17] = 8'd197;
	sample_rom[75][18] = 8'd219;
	sample_rom[75][19] = 8'd231;
	sample_rom[75][20] = 8'd235;
	sample_rom[75][21] = 8'd231;
	sample_rom[75][22] = 8'd219;
	sample_rom[75][23] = 8'd201;
	sample_rom[75][24] = 8'd179;
	sample_rom[75][25] = 8'd159;
	sample_rom[75][26] = 8'd140;
	sample_rom[75][27] = 8'd131;
	sample_rom[75][28] = 8'd126;
	sample_rom[75][29] = 8'd133;
	sample_rom[75][30] = 8'd146;
	sample_rom[75][31] = 8'd163;
	sample_rom[75][32] = 8'd186;
	sample_rom[75][33] = 8'd207;
	sample_rom[75][34] = 8'd225;
	sample_rom[75][35] = 8'd235;
	sample_rom[75][36] = 8'd239;
	sample_rom[75][37] = 8'd233;
	sample_rom[75][38] = 8'd221;
	sample_rom[75][39] = 8'd200;
	sample_rom[75][40] = 8'd179;
	sample_rom[75][41] = 8'd156;
	sample_rom[75][42] = 8'd138;
	sample_rom[75][43] = 8'd125;
	sample_rom[75][44] = 8'd120;
	sample_rom[75][45] = 8'd126;
	sample_rom[75][46] = 8'd138;
	sample_rom[75][47] = 8'd153;
	sample_rom[75][48] = 8'd170;
	sample_rom[75][49] = 8'd189;
	sample_rom[75][50] = 8'd202;
	sample_rom[75][51] = 8'd207;
	sample_rom[75][52] = 8'd208;
	sample_rom[75][53] = 8'd200;
	sample_rom[75][54] = 8'd186;
	sample_rom[75][55] = 8'd165;
	sample_rom[75][56] = 8'd146;
	sample_rom[75][57] = 8'd125;
	sample_rom[75][58] = 8'd107;
	sample_rom[75][59] = 8'd98;
	sample_rom[75][60] = 8'd93;
	sample_rom[75][61] = 8'd96;
	sample_rom[75][62] = 8'd100;
	sample_rom[75][63] = 8'd112;
	sample_rom[76][0] = 8'd130;
	sample_rom[76][1] = 8'd163;
	sample_rom[76][2] = 8'd191;
	sample_rom[76][3] = 8'd206;
	sample_rom[76][4] = 8'd208;
	sample_rom[76][5] = 8'd196;
	sample_rom[76][6] = 8'd174;
	sample_rom[76][7] = 8'd148;
	sample_rom[76][8] = 8'd121;
	sample_rom[76][9] = 8'd101;
	sample_rom[76][10] = 8'd93;
	sample_rom[76][11] = 8'd94;
	sample_rom[76][12] = 8'd108;
	sample_rom[76][13] = 8'd134;
	sample_rom[76][14] = 8'd163;
	sample_rom[76][15] = 8'd193;
	sample_rom[76][16] = 8'd218;
	sample_rom[76][17] = 8'd231;
	sample_rom[76][18] = 8'd232;
	sample_rom[76][19] = 8'd224;
	sample_rom[76][20] = 8'd207;
	sample_rom[76][21] = 8'd183;
	sample_rom[76][22] = 8'd159;
	sample_rom[76][23] = 8'd139;
	sample_rom[76][24] = 8'd126;
	sample_rom[76][25] = 8'd125;
	sample_rom[76][26] = 8'd134;
	sample_rom[76][27] = 8'd152;
	sample_rom[76][28] = 8'd174;
	sample_rom[76][29] = 8'd200;
	sample_rom[76][30] = 8'd222;
	sample_rom[76][31] = 8'd235;
	sample_rom[76][32] = 8'd240;
	sample_rom[76][33] = 8'd232;
	sample_rom[76][34] = 8'd218;
	sample_rom[76][35] = 8'd196;
	sample_rom[76][36] = 8'd170;
	sample_rom[76][37] = 8'd149;
	sample_rom[76][38] = 8'd136;
	sample_rom[76][39] = 8'd127;
	sample_rom[76][40] = 8'd134;
	sample_rom[76][41] = 8'd145;
	sample_rom[76][42] = 8'd166;
	sample_rom[76][43] = 8'd186;
	sample_rom[76][44] = 8'd204;
	sample_rom[76][45] = 8'd216;
	sample_rom[76][46] = 8'd221;
	sample_rom[76][47] = 8'd213;
	sample_rom[76][48] = 8'd198;
	sample_rom[76][49] = 8'd176;
	sample_rom[76][50] = 8'd155;
	sample_rom[76][51] = 8'd133;
	sample_rom[76][52] = 8'd120;
	sample_rom[76][53] = 8'd113;
	sample_rom[76][54] = 8'd114;
	sample_rom[76][55] = 8'd121;
	sample_rom[76][56] = 8'd136;
	sample_rom[76][57] = 8'd152;
	sample_rom[76][58] = 8'd165;
	sample_rom[76][59] = 8'd175;
	sample_rom[76][60] = 8'd178;
	sample_rom[76][61] = 8'd173;
	sample_rom[76][62] = 8'd162;
	sample_rom[76][63] = 8'd145;
	sample_rom[77][0] = 8'd130;
	sample_rom[77][1] = 8'd142;
	sample_rom[77][2] = 8'd153;
	sample_rom[77][3] = 8'd160;
	sample_rom[77][4] = 8'd164;
	sample_rom[77][5] = 8'd164;
	sample_rom[77][6] = 8'd164;
	sample_rom[77][7] = 8'd161;
	sample_rom[77][8] = 8'd160;
	sample_rom[77][9] = 8'd159;
	sample_rom[77][10] = 8'd160;
	sample_rom[77][11] = 8'd164;
	sample_rom[77][12] = 8'd170;
	sample_rom[77][13] = 8'd178;
	sample_rom[77][14] = 8'd189;
	sample_rom[77][15] = 8'd200;
	sample_rom[77][16] = 8'd208;
	sample_rom[77][17] = 8'd215;
	sample_rom[77][18] = 8'd217;
	sample_rom[77][19] = 8'd218;
	sample_rom[77][20] = 8'd215;
	sample_rom[77][21] = 8'd213;
	sample_rom[77][22] = 8'd207;
	sample_rom[77][23] = 8'd204;
	sample_rom[77][24] = 8'd202;
	sample_rom[77][25] = 8'd203;
	sample_rom[77][26] = 8'd206;
	sample_rom[77][27] = 8'd212;
	sample_rom[77][28] = 8'd219;
	sample_rom[77][29] = 8'd225;
	sample_rom[77][30] = 8'd232;
	sample_rom[77][31] = 8'd236;
	sample_rom[77][32] = 8'd237;
	sample_rom[77][33] = 8'd236;
	sample_rom[77][34] = 8'd231;
	sample_rom[77][35] = 8'd225;
	sample_rom[77][36] = 8'd218;
	sample_rom[77][37] = 8'd210;
	sample_rom[77][38] = 8'd204;
	sample_rom[77][39] = 8'd201;
	sample_rom[77][40] = 8'd201;
	sample_rom[77][41] = 8'd202;
	sample_rom[77][42] = 8'd207;
	sample_rom[77][43] = 8'd210;
	sample_rom[77][44] = 8'd214;
	sample_rom[77][45] = 8'd215;
	sample_rom[77][46] = 8'd215;
	sample_rom[77][47] = 8'd211;
	sample_rom[77][48] = 8'd205;
	sample_rom[77][49] = 8'd195;
	sample_rom[77][50] = 8'd184;
	sample_rom[77][51] = 8'd174;
	sample_rom[77][52] = 8'd166;
	sample_rom[77][53] = 8'd160;
	sample_rom[77][54] = 8'd156;
	sample_rom[77][55] = 8'd155;
	sample_rom[77][56] = 8'd157;
	sample_rom[77][57] = 8'd159;
	sample_rom[77][58] = 8'd160;
	sample_rom[77][59] = 8'd162;
	sample_rom[77][60] = 8'd160;
	sample_rom[77][61] = 8'd156;
	sample_rom[77][62] = 8'd147;
	sample_rom[77][63] = 8'd136;
	sample_rom[78][0] = 8'd130;
	sample_rom[78][1] = 8'd146;
	sample_rom[78][2] = 8'd158;
	sample_rom[78][3] = 8'd167;
	sample_rom[78][4] = 8'd174;
	sample_rom[78][5] = 8'd178;
	sample_rom[78][6] = 8'd179;
	sample_rom[78][7] = 8'd179;
	sample_rom[78][8] = 8'd178;
	sample_rom[78][9] = 8'd177;
	sample_rom[78][10] = 8'd179;
	sample_rom[78][11] = 8'd184;
	sample_rom[78][12] = 8'd190;
	sample_rom[78][13] = 8'd198;
	sample_rom[78][14] = 8'd208;
	sample_rom[78][15] = 8'd218;
	sample_rom[78][16] = 8'd223;
	sample_rom[78][17] = 8'd227;
	sample_rom[78][18] = 8'd227;
	sample_rom[78][19] = 8'd225;
	sample_rom[78][20] = 8'd220;
	sample_rom[78][21] = 8'd212;
	sample_rom[78][22] = 8'd203;
	sample_rom[78][23] = 8'd195;
	sample_rom[78][24] = 8'd189;
	sample_rom[78][25] = 8'd185;
	sample_rom[78][26] = 8'd182;
	sample_rom[78][27] = 8'd182;
	sample_rom[78][28] = 8'd183;
	sample_rom[78][29] = 8'd184;
	sample_rom[78][30] = 8'd185;
	sample_rom[78][31] = 8'd183;
	sample_rom[78][32] = 8'd179;
	sample_rom[78][33] = 8'd172;
	sample_rom[78][34] = 8'd162;
	sample_rom[78][35] = 8'd152;
	sample_rom[78][36] = 8'd140;
	sample_rom[78][37] = 8'd127;
	sample_rom[78][38] = 8'd118;
	sample_rom[78][39] = 8'd111;
	sample_rom[78][40] = 8'd107;
	sample_rom[78][41] = 8'd107;
	sample_rom[78][42] = 8'd109;
	sample_rom[78][43] = 8'd112;
	sample_rom[78][44] = 8'd115;
	sample_rom[78][45] = 8'd116;
	sample_rom[78][46] = 8'd115;
	sample_rom[78][47] = 8'd112;
	sample_rom[78][48] = 8'd108;
	sample_rom[78][49] = 8'd101;
	sample_rom[78][50] = 8'd95;
	sample_rom[78][51] = 8'd88;
	sample_rom[78][52] = 8'd85;
	sample_rom[78][53] = 8'd83;
	sample_rom[78][54] = 8'd84;
	sample_rom[78][55] = 8'd89;
	sample_rom[78][56] = 8'd97;
	sample_rom[78][57] = 8'd105;
	sample_rom[78][58] = 8'd115;
	sample_rom[78][59] = 8'd124;
	sample_rom[78][60] = 8'd129;
	sample_rom[78][61] = 8'd133;
	sample_rom[78][62] = 8'd133;
	sample_rom[78][63] = 8'd131;
	sample_rom[79][0] = 8'd130;
	sample_rom[79][1] = 8'd149;
	sample_rom[79][2] = 8'd163;
	sample_rom[79][3] = 8'd175;
	sample_rom[79][4] = 8'd183;
	sample_rom[79][5] = 8'd187;
	sample_rom[79][6] = 8'd187;
	sample_rom[79][7] = 8'd186;
	sample_rom[79][8] = 8'd184;
	sample_rom[79][9] = 8'd185;
	sample_rom[79][10] = 8'd189;
	sample_rom[79][11] = 8'd194;
	sample_rom[79][12] = 8'd200;
	sample_rom[79][13] = 8'd206;
	sample_rom[79][14] = 8'd211;
	sample_rom[79][15] = 8'd213;
	sample_rom[79][16] = 8'd210;
	sample_rom[79][17] = 8'd202;
	sample_rom[79][18] = 8'd191;
	sample_rom[79][19] = 8'd177;
	sample_rom[79][20] = 8'd163;
	sample_rom[79][21] = 8'd150;
	sample_rom[79][22] = 8'd140;
	sample_rom[79][23] = 8'd133;
	sample_rom[79][24] = 8'd130;
	sample_rom[79][25] = 8'd130;
	sample_rom[79][26] = 8'd131;
	sample_rom[79][27] = 8'd132;
	sample_rom[79][28] = 8'd132;
	sample_rom[79][29] = 8'd129;
	sample_rom[79][30] = 8'd124;
	sample_rom[79][31] = 8'd116;
	sample_rom[79][32] = 8'd108;
	sample_rom[79][33] = 8'd101;
	sample_rom[79][34] = 8'd98;
	sample_rom[79][35] = 8'd100;
	sample_rom[79][36] = 8'd105;
	sample_rom[79][37] = 8'd114;
	sample_rom[79][38] = 8'd126;
	sample_rom[79][39] = 8'd140;
	sample_rom[79][40] = 8'd153;
	sample_rom[79][41] = 8'd163;
	sample_rom[79][42] = 8'd171;
	sample_rom[79][43] = 8'd175;
	sample_rom[79][44] = 8'd177;
	sample_rom[79][45] = 8'd176;
	sample_rom[79][46] = 8'd176;
	sample_rom[79][47] = 8'd177;
	sample_rom[79][48] = 8'd181;
	sample_rom[79][49] = 8'd186;
	sample_rom[79][50] = 8'd194;
	sample_rom[79][51] = 8'd203;
	sample_rom[79][52] = 8'd211;
	sample_rom[79][53] = 8'd216;
	sample_rom[79][54] = 8'd216;
	sample_rom[79][55] = 8'd212;
	sample_rom[79][56] = 8'd205;
	sample_rom[79][57] = 8'd191;
	sample_rom[79][58] = 8'd178;
	sample_rom[79][59] = 8'd164;
	sample_rom[79][60] = 8'd152;
	sample_rom[79][61] = 8'd141;
	sample_rom[79][62] = 8'd134;
	sample_rom[79][63] = 8'd130;
	sample_rom[80][0] = 8'd130;
	sample_rom[80][1] = 8'd148;
	sample_rom[80][2] = 8'd161;
	sample_rom[80][3] = 8'd174;
	sample_rom[80][4] = 8'd179;
	sample_rom[80][5] = 8'd180;
	sample_rom[80][6] = 8'd179;
	sample_rom[80][7] = 8'd178;
	sample_rom[80][8] = 8'd176;
	sample_rom[80][9] = 8'd175;
	sample_rom[80][10] = 8'd178;
	sample_rom[80][11] = 8'd179;
	sample_rom[80][12] = 8'd181;
	sample_rom[80][13] = 8'd181;
	sample_rom[80][14] = 8'd177;
	sample_rom[80][15] = 8'd169;
	sample_rom[80][16] = 8'd159;
	sample_rom[80][17] = 8'd144;
	sample_rom[80][18] = 8'd130;
	sample_rom[80][19] = 8'd118;
	sample_rom[80][20] = 8'd108;
	sample_rom[80][21] = 8'd104;
	sample_rom[80][22] = 8'd104;
	sample_rom[80][23] = 8'd108;
	sample_rom[80][24] = 8'd114;
	sample_rom[80][25] = 8'd122;
	sample_rom[80][26] = 8'd128;
	sample_rom[80][27] = 8'd131;
	sample_rom[80][28] = 8'd133;
	sample_rom[80][29] = 8'd135;
	sample_rom[80][30] = 8'd137;
	sample_rom[80][31] = 8'd141;
	sample_rom[80][32] = 8'd148;
	sample_rom[80][33] = 8'd160;
	sample_rom[80][34] = 8'd172;
	sample_rom[80][35] = 8'd187;
	sample_rom[80][36] = 8'd200;
	sample_rom[80][37] = 8'd210;
	sample_rom[80][38] = 8'd214;
	sample_rom[80][39] = 8'd213;
	sample_rom[80][40] = 8'd209;
	sample_rom[80][41] = 8'd199;
	sample_rom[80][42] = 8'd191;
	sample_rom[80][43] = 8'd181;
	sample_rom[80][44] = 8'd174;
	sample_rom[80][45] = 8'd168;
	sample_rom[80][46] = 8'd165;
	sample_rom[80][47] = 8'd161;
	sample_rom[80][48] = 8'd158;
	sample_rom[80][49] = 8'd150;
	sample_rom[80][50] = 8'd141;
	sample_rom[80][51] = 8'd127;
	sample_rom[80][52] = 8'd112;
	sample_rom[80][53] = 8'd99;
	sample_rom[80][54] = 8'd89;
	sample_rom[80][55] = 8'd82;
	sample_rom[80][56] = 8'd81;
	sample_rom[80][57] = 8'd86;
	sample_rom[80][58] = 8'd92;
	sample_rom[80][59] = 8'd102;
	sample_rom[80][60] = 8'd112;
	sample_rom[80][61] = 8'd120;
	sample_rom[80][62] = 8'd124;
	sample_rom[80][63] = 8'd127;
	sample_rom[81][0] = 8'd130;
	sample_rom[81][1] = 8'd155;
	sample_rom[81][2] = 8'd175;
	sample_rom[81][3] = 8'd189;
	sample_rom[81][4] = 8'd195;
	sample_rom[81][5] = 8'd195;
	sample_rom[81][6] = 8'd191;
	sample_rom[81][7] = 8'd185;
	sample_rom[81][8] = 8'd180;
	sample_rom[81][9] = 8'd177;
	sample_rom[81][10] = 8'd177;
	sample_rom[81][11] = 8'd175;
	sample_rom[81][12] = 8'd170;
	sample_rom[81][13] = 8'd162;
	sample_rom[81][14] = 8'd149;
	sample_rom[81][15] = 8'd132;
	sample_rom[81][16] = 8'd114;
	sample_rom[81][17] = 8'd98;
	sample_rom[81][18] = 8'd90;
	sample_rom[81][19] = 8'd87;
	sample_rom[81][20] = 8'd94;
	sample_rom[81][21] = 8'd107;
	sample_rom[81][22] = 8'd124;
	sample_rom[81][23] = 8'd143;
	sample_rom[81][24] = 8'd158;
	sample_rom[81][25] = 8'd170;
	sample_rom[81][26] = 8'd178;
	sample_rom[81][27] = 8'd183;
	sample_rom[81][28] = 8'd187;
	sample_rom[81][29] = 8'd194;
	sample_rom[81][30] = 8'd202;
	sample_rom[81][31] = 8'd213;
	sample_rom[81][32] = 8'd223;
	sample_rom[81][33] = 8'd228;
	sample_rom[81][34] = 8'd228;
	sample_rom[81][35] = 8'd222;
	sample_rom[81][36] = 8'd207;
	sample_rom[81][37] = 8'd185;
	sample_rom[81][38] = 8'd162;
	sample_rom[81][39] = 8'd141;
	sample_rom[81][40] = 8'd125;
	sample_rom[81][41] = 8'd114;
	sample_rom[81][42] = 8'd111;
	sample_rom[81][43] = 8'd112;
	sample_rom[81][44] = 8'd113;
	sample_rom[81][45] = 8'd115;
	sample_rom[81][46] = 8'd116;
	sample_rom[81][47] = 8'd116;
	sample_rom[81][48] = 8'd115;
	sample_rom[81][49] = 8'd115;
	sample_rom[81][50] = 8'd123;
	sample_rom[81][51] = 8'd134;
	sample_rom[81][52] = 8'd151;
	sample_rom[81][53] = 8'd169;
	sample_rom[81][54] = 8'd188;
	sample_rom[81][55] = 8'd202;
	sample_rom[81][56] = 8'd209;
	sample_rom[81][57] = 8'd209;
	sample_rom[81][58] = 8'd200;
	sample_rom[81][59] = 8'd186;
	sample_rom[81][60] = 8'd170;
	sample_rom[81][61] = 8'd156;
	sample_rom[81][62] = 8'd143;
	sample_rom[81][63] = 8'd134;
	sample_rom[82][0] = 8'd130;
	sample_rom[82][1] = 8'd159;
	sample_rom[82][2] = 8'd180;
	sample_rom[82][3] = 8'd193;
	sample_rom[82][4] = 8'd197;
	sample_rom[82][5] = 8'd194;
	sample_rom[82][6] = 8'd185;
	sample_rom[82][7] = 8'd176;
	sample_rom[82][8] = 8'd168;
	sample_rom[82][9] = 8'd162;
	sample_rom[82][10] = 8'd159;
	sample_rom[82][11] = 8'd153;
	sample_rom[82][12] = 8'd142;
	sample_rom[82][13] = 8'd128;
	sample_rom[82][14] = 8'd112;
	sample_rom[82][15] = 8'd97;
	sample_rom[82][16] = 8'd88;
	sample_rom[82][17] = 8'd88;
	sample_rom[82][18] = 8'd98;
	sample_rom[82][19] = 8'd117;
	sample_rom[82][20] = 8'd143;
	sample_rom[82][21] = 8'd168;
	sample_rom[82][22] = 8'd189;
	sample_rom[82][23] = 8'd204;
	sample_rom[82][24] = 8'd211;
	sample_rom[82][25] = 8'd211;
	sample_rom[82][26] = 8'd209;
	sample_rom[82][27] = 8'd207;
	sample_rom[82][28] = 8'd206;
	sample_rom[82][29] = 8'd204;
	sample_rom[82][30] = 8'd201;
	sample_rom[82][31] = 8'd193;
	sample_rom[82][32] = 8'd179;
	sample_rom[82][33] = 8'd160;
	sample_rom[82][34] = 8'd137;
	sample_rom[82][35] = 8'd116;
	sample_rom[82][36] = 8'd100;
	sample_rom[82][37] = 8'd93;
	sample_rom[82][38] = 8'd97;
	sample_rom[82][39] = 8'd111;
	sample_rom[82][40] = 8'd129;
	sample_rom[82][41] = 8'd149;
	sample_rom[82][42] = 8'd165;
	sample_rom[82][43] = 8'd178;
	sample_rom[82][44] = 8'd184;
	sample_rom[82][45] = 8'd188;
	sample_rom[82][46] = 8'd190;
	sample_rom[82][47] = 8'd195;
	sample_rom[82][48] = 8'd201;
	sample_rom[82][49] = 8'd205;
	sample_rom[82][50] = 8'd206;
	sample_rom[82][51] = 8'd199;
	sample_rom[82][52] = 8'd184;
	sample_rom[82][53] = 8'd160;
	sample_rom[82][54] = 8'd133;
	sample_rom[82][55] = 8'd106;
	sample_rom[82][56] = 8'd87;
	sample_rom[82][57] = 8'd75;
	sample_rom[82][58] = 8'd73;
	sample_rom[82][59] = 8'd81;
	sample_rom[82][60] = 8'd93;
	sample_rom[82][61] = 8'd104;
	sample_rom[82][62] = 8'd115;
	sample_rom[82][63] = 8'd123;
	sample_rom[83][0] = 8'd130;
	sample_rom[83][1] = 8'd161;
	sample_rom[83][2] = 8'd185;
	sample_rom[83][3] = 8'd197;
	sample_rom[83][4] = 8'd199;
	sample_rom[83][5] = 8'd189;
	sample_rom[83][6] = 8'd176;
	sample_rom[83][7] = 8'd164;
	sample_rom[83][8] = 8'd153;
	sample_rom[83][9] = 8'd145;
	sample_rom[83][10] = 8'd138;
	sample_rom[83][11] = 8'd128;
	sample_rom[83][12] = 8'd116;
	sample_rom[83][13] = 8'd103;
	sample_rom[83][14] = 8'd94;
	sample_rom[83][15] = 8'd93;
	sample_rom[83][16] = 8'd101;
	sample_rom[83][17] = 8'd122;
	sample_rom[83][18] = 8'd151;
	sample_rom[83][19] = 8'd181;
	sample_rom[83][20] = 8'd206;
	sample_rom[83][21] = 8'd222;
	sample_rom[83][22] = 8'd223;
	sample_rom[83][23] = 8'd218;
	sample_rom[83][24] = 8'd205;
	sample_rom[83][25] = 8'd191;
	sample_rom[83][26] = 8'd178;
	sample_rom[83][27] = 8'd169;
	sample_rom[83][28] = 8'd159;
	sample_rom[83][29] = 8'd149;
	sample_rom[83][30] = 8'd136;
	sample_rom[83][31] = 8'd121;
	sample_rom[83][32] = 8'd108;
	sample_rom[83][33] = 8'd103;
	sample_rom[83][34] = 8'd107;
	sample_rom[83][35] = 8'd124;
	sample_rom[83][36] = 8'd151;
	sample_rom[83][37] = 8'd179;
	sample_rom[83][38] = 8'd206;
	sample_rom[83][39] = 8'd222;
	sample_rom[83][40] = 8'd225;
	sample_rom[83][41] = 8'd220;
	sample_rom[83][42] = 8'd206;
	sample_rom[83][43] = 8'd189;
	sample_rom[83][44] = 8'd175;
	sample_rom[83][45] = 8'd163;
	sample_rom[83][46] = 8'd154;
	sample_rom[83][47] = 8'd142;
	sample_rom[83][48] = 8'd128;
	sample_rom[83][49] = 8'd113;
	sample_rom[83][50] = 8'd97;
	sample_rom[83][51] = 8'd88;
	sample_rom[83][52] = 8'd89;
	sample_rom[83][53] = 8'd99;
	sample_rom[83][54] = 8'd122;
	sample_rom[83][55] = 8'd149;
	sample_rom[83][56] = 8'd175;
	sample_rom[83][57] = 8'd194;
	sample_rom[83][58] = 8'd201;
	sample_rom[83][59] = 8'd197;
	sample_rom[83][60] = 8'd184;
	sample_rom[83][61] = 8'd166;
	sample_rom[83][62] = 8'd152;
	sample_rom[83][63] = 8'd138;
	sample_rom[84][0] = 8'd130;
	sample_rom[84][1] = 8'd158;
	sample_rom[84][2] = 8'd179;
	sample_rom[84][3] = 8'd187;
	sample_rom[84][4] = 8'd184;
	sample_rom[84][5] = 8'd172;
	sample_rom[84][6] = 8'd159;
	sample_rom[84][7] = 8'd146;
	sample_rom[84][8] = 8'd135;
	sample_rom[84][9] = 8'd128;
	sample_rom[84][10] = 8'd120;
	sample_rom[84][11] = 8'd113;
	sample_rom[84][12] = 8'd105;
	sample_rom[84][13] = 8'd102;
	sample_rom[84][14] = 8'd106;
	sample_rom[84][15] = 8'd120;
	sample_rom[84][16] = 8'd143;
	sample_rom[84][17] = 8'd170;
	sample_rom[84][18] = 8'd195;
	sample_rom[84][19] = 8'd210;
	sample_rom[84][20] = 8'd212;
	sample_rom[84][21] = 8'd202;
	sample_rom[84][22] = 8'd182;
	sample_rom[84][23] = 8'd161;
	sample_rom[84][24] = 8'd144;
	sample_rom[84][25] = 8'd134;
	sample_rom[84][26] = 8'd128;
	sample_rom[84][27] = 8'd126;
	sample_rom[84][28] = 8'd123;
	sample_rom[84][29] = 8'd123;
	sample_rom[84][30] = 8'd125;
	sample_rom[84][31] = 8'd134;
	sample_rom[84][32] = 8'd148;
	sample_rom[84][33] = 8'd169;
	sample_rom[84][34] = 8'd193;
	sample_rom[84][35] = 8'd210;
	sample_rom[84][36] = 8'd219;
	sample_rom[84][37] = 8'd213;
	sample_rom[84][38] = 8'd193;
	sample_rom[84][39] = 8'd167;
	sample_rom[84][40] = 8'd144;
	sample_rom[84][41] = 8'd125;
	sample_rom[84][42] = 8'd115;
	sample_rom[84][43] = 8'd114;
	sample_rom[84][44] = 8'd117;
	sample_rom[84][45] = 8'd122;
	sample_rom[84][46] = 8'd127;
	sample_rom[84][47] = 8'd133;
	sample_rom[84][48] = 8'd142;
	sample_rom[84][49] = 8'd155;
	sample_rom[84][50] = 8'd173;
	sample_rom[84][51] = 8'd187;
	sample_rom[84][52] = 8'd199;
	sample_rom[84][53] = 8'd199;
	sample_rom[84][54] = 8'd185;
	sample_rom[84][55] = 8'd161;
	sample_rom[84][56] = 8'd134;
	sample_rom[84][57] = 8'd107;
	sample_rom[84][58] = 8'd90;
	sample_rom[84][59] = 8'd86;
	sample_rom[84][60] = 8'd90;
	sample_rom[84][61] = 8'd98;
	sample_rom[84][62] = 8'd110;
	sample_rom[84][63] = 8'd120;
	sample_rom[85][0] = 8'd135;
	sample_rom[85][1] = 8'd184;
	sample_rom[85][2] = 8'd218;
	sample_rom[85][3] = 8'd228;
	sample_rom[85][4] = 8'd219;
	sample_rom[85][5] = 8'd197;
	sample_rom[85][6] = 8'd180;
	sample_rom[85][7] = 8'd176;
	sample_rom[85][8] = 8'd183;
	sample_rom[85][9] = 8'd196;
	sample_rom[85][10] = 8'd206;
	sample_rom[85][11] = 8'd207;
	sample_rom[85][12] = 8'd199;
	sample_rom[85][13] = 8'd189;
	sample_rom[85][14] = 8'd181;
	sample_rom[85][15] = 8'd184;
	sample_rom[85][16] = 8'd193;
	sample_rom[85][17] = 8'd201;
	sample_rom[85][18] = 8'd199;
	sample_rom[85][19] = 8'd189;
	sample_rom[85][20] = 8'd173;
	sample_rom[85][21] = 8'd160;
	sample_rom[85][22] = 8'd155;
	sample_rom[85][23] = 8'd157;
	sample_rom[85][24] = 8'd160;
	sample_rom[85][25] = 8'd160;
	sample_rom[85][26] = 8'd140;
	sample_rom[85][27] = 8'd113;
	sample_rom[85][28] = 8'd81;
	sample_rom[85][29] = 8'd63;
	sample_rom[85][30] = 8'd64;
	sample_rom[85][31] = 8'd89;
	sample_rom[85][32] = 8'd131;
	sample_rom[85][33] = 8'd171;
	sample_rom[85][34] = 8'd195;
	sample_rom[85][35] = 8'd198;
	sample_rom[85][36] = 8'd179;
	sample_rom[85][37] = 8'd152;
	sample_rom[85][38] = 8'd129;
	sample_rom[85][39] = 8'd120;
	sample_rom[85][40] = 8'd123;
	sample_rom[85][41] = 8'd135;
	sample_rom[85][42] = 8'd142;
	sample_rom[85][43] = 8'd144;
	sample_rom[85][44] = 8'd136;
	sample_rom[85][45] = 8'd127;
	sample_rom[85][46] = 8'd123;
	sample_rom[85][47] = 8'd128;
	sample_rom[85][48] = 8'd140;
	sample_rom[85][49] = 8'd151;
	sample_rom[85][50] = 8'd156;
	sample_rom[85][51] = 8'd150;
	sample_rom[85][52] = 8'd137;
	sample_rom[85][53] = 8'd130;
	sample_rom[85][54] = 8'd129;
	sample_rom[85][55] = 8'd135;
	sample_rom[85][56] = 8'd144;
	sample_rom[85][57] = 8'd145;
	sample_rom[85][58] = 8'd132;
	sample_rom[85][59] = 8'd107;
	sample_rom[85][60] = 8'd77;
	sample_rom[85][61] = 8'd61;
	sample_rom[85][62] = 8'd62;
	sample_rom[85][63] = 8'd90;
	sample_rom[86][0] = 8'd132;
	sample_rom[86][1] = 8'd169;
	sample_rom[86][2] = 8'd200;
	sample_rom[86][3] = 8'd224;
	sample_rom[86][4] = 8'd239;
	sample_rom[86][5] = 8'd246;
	sample_rom[86][6] = 8'd247;
	sample_rom[86][7] = 8'd243;
	sample_rom[86][8] = 8'd236;
	sample_rom[86][9] = 8'd231;
	sample_rom[86][10] = 8'd226;
	sample_rom[86][11] = 8'd223;
	sample_rom[86][12] = 8'd221;
	sample_rom[86][13] = 8'd220;
	sample_rom[86][14] = 8'd221;
	sample_rom[86][15] = 8'd218;
	sample_rom[86][16] = 8'd217;
	sample_rom[86][17] = 8'd215;
	sample_rom[86][18] = 8'd212;
	sample_rom[86][19] = 8'd205;
	sample_rom[86][20] = 8'd202;
	sample_rom[86][21] = 8'd193;
	sample_rom[86][22] = 8'd189;
	sample_rom[86][23] = 8'd185;
	sample_rom[86][24] = 8'd182;
	sample_rom[86][25] = 8'd177;
	sample_rom[86][26] = 8'd173;
	sample_rom[86][27] = 8'd172;
	sample_rom[86][28] = 8'd166;
	sample_rom[86][29] = 8'd162;
	sample_rom[86][30] = 8'd159;
	sample_rom[86][31] = 8'd155;
	sample_rom[86][32] = 8'd155;
	sample_rom[86][33] = 8'd157;
	sample_rom[86][34] = 8'd159;
	sample_rom[86][35] = 8'd160;
	sample_rom[86][36] = 8'd164;
	sample_rom[86][37] = 8'd163;
	sample_rom[86][38] = 8'd163;
	sample_rom[86][39] = 8'd160;
	sample_rom[86][40] = 8'd159;
	sample_rom[86][41] = 8'd156;
	sample_rom[86][42] = 8'd155;
	sample_rom[86][43] = 8'd153;
	sample_rom[86][44] = 8'd150;
	sample_rom[86][45] = 8'd150;
	sample_rom[86][46] = 8'd147;
	sample_rom[86][47] = 8'd141;
	sample_rom[86][48] = 8'd137;
	sample_rom[86][49] = 8'd132;
	sample_rom[86][50] = 8'd129;
	sample_rom[86][51] = 8'd129;
	sample_rom[86][52] = 8'd128;
	sample_rom[86][53] = 8'd127;
	sample_rom[86][54] = 8'd126;
	sample_rom[86][55] = 8'd125;
	sample_rom[86][56] = 8'd124;
	sample_rom[86][57] = 8'd124;
	sample_rom[86][58] = 8'd124;
	sample_rom[86][59] = 8'd127;
	sample_rom[86][60] = 8'd127;
	sample_rom[86][61] = 8'd131;
	sample_rom[86][62] = 8'd128;
	sample_rom[86][63] = 8'd129;
	sample_rom[87][0] = 8'd132;
	sample_rom[87][1] = 8'd167;
	sample_rom[87][2] = 8'd197;
	sample_rom[87][3] = 8'd220;
	sample_rom[87][4] = 8'd230;
	sample_rom[87][5] = 8'd236;
	sample_rom[87][6] = 8'd232;
	sample_rom[87][7] = 8'd223;
	sample_rom[87][8] = 8'd213;
	sample_rom[87][9] = 8'd203;
	sample_rom[87][10] = 8'd195;
	sample_rom[87][11] = 8'd190;
	sample_rom[87][12] = 8'd190;
	sample_rom[87][13] = 8'd186;
	sample_rom[87][14] = 8'd189;
	sample_rom[87][15] = 8'd186;
	sample_rom[87][16] = 8'd182;
	sample_rom[87][17] = 8'd178;
	sample_rom[87][18] = 8'd174;
	sample_rom[87][19] = 8'd166;
	sample_rom[87][20] = 8'd164;
	sample_rom[87][21] = 8'd160;
	sample_rom[87][22] = 8'd159;
	sample_rom[87][23] = 8'd158;
	sample_rom[87][24] = 8'd156;
	sample_rom[87][25] = 8'd153;
	sample_rom[87][26] = 8'd146;
	sample_rom[87][27] = 8'd140;
	sample_rom[87][28] = 8'd130;
	sample_rom[87][29] = 8'd125;
	sample_rom[87][30] = 8'd121;
	sample_rom[87][31] = 8'd119;
	sample_rom[87][32] = 8'd120;
	sample_rom[87][33] = 8'd122;
	sample_rom[87][34] = 8'd128;
	sample_rom[87][35] = 8'd132;
	sample_rom[87][36] = 8'd140;
	sample_rom[87][37] = 8'd141;
	sample_rom[87][38] = 8'd143;
	sample_rom[87][39] = 8'd143;
	sample_rom[87][40] = 8'd144;
	sample_rom[87][41] = 8'd144;
	sample_rom[87][42] = 8'd144;
	sample_rom[87][43] = 8'd143;
	sample_rom[87][44] = 8'd145;
	sample_rom[87][45] = 8'd143;
	sample_rom[87][46] = 8'd138;
	sample_rom[87][47] = 8'd136;
	sample_rom[87][48] = 8'd130;
	sample_rom[87][49] = 8'd125;
	sample_rom[87][50] = 8'd122;
	sample_rom[87][51] = 8'd116;
	sample_rom[87][52] = 8'd115;
	sample_rom[87][53] = 8'd115;
	sample_rom[87][54] = 8'd117;
	sample_rom[87][55] = 8'd119;
	sample_rom[87][56] = 8'd123;
	sample_rom[87][57] = 8'd124;
	sample_rom[87][58] = 8'd126;
	sample_rom[87][59] = 8'd131;
	sample_rom[87][60] = 8'd132;
	sample_rom[87][61] = 8'd131;
	sample_rom[87][62] = 8'd131;
	sample_rom[87][63] = 8'd131;
	sample_rom[88][0] = 8'd131;
	sample_rom[88][1] = 8'd168;
	sample_rom[88][2] = 8'd199;
	sample_rom[88][3] = 8'd217;
	sample_rom[88][4] = 8'd223;
	sample_rom[88][5] = 8'd223;
	sample_rom[88][6] = 8'd218;
	sample_rom[88][7] = 8'd217;
	sample_rom[88][8] = 8'd219;
	sample_rom[88][9] = 8'd223;
	sample_rom[88][10] = 8'd228;
	sample_rom[88][11] = 8'd231;
	sample_rom[88][12] = 8'd235;
	sample_rom[88][13] = 8'd235;
	sample_rom[88][14] = 8'd232;
	sample_rom[88][15] = 8'd232;
	sample_rom[88][16] = 8'd224;
	sample_rom[88][17] = 8'd223;
	sample_rom[88][18] = 8'd217;
	sample_rom[88][19] = 8'd212;
	sample_rom[88][20] = 8'd212;
	sample_rom[88][21] = 8'd209;
	sample_rom[88][22] = 8'd211;
	sample_rom[88][23] = 8'd216;
	sample_rom[88][24] = 8'd214;
	sample_rom[88][25] = 8'd214;
	sample_rom[88][26] = 8'd212;
	sample_rom[88][27] = 8'd210;
	sample_rom[88][28] = 8'd210;
	sample_rom[88][29] = 8'd207;
	sample_rom[88][30] = 8'd207;
	sample_rom[88][31] = 8'd204;
	sample_rom[88][32] = 8'd202;
	sample_rom[88][33] = 8'd195;
	sample_rom[88][34] = 8'd188;
	sample_rom[88][35] = 8'd181;
	sample_rom[88][36] = 8'd173;
	sample_rom[88][37] = 8'd173;
	sample_rom[88][38] = 8'd175;
	sample_rom[88][39] = 8'd175;
	sample_rom[88][40] = 8'd176;
	sample_rom[88][41] = 8'd178;
	sample_rom[88][42] = 8'd178;
	sample_rom[88][43] = 8'd173;
	sample_rom[88][44] = 8'd173;
	sample_rom[88][45] = 8'd171;
	sample_rom[88][46] = 8'd166;
	sample_rom[88][47] = 8'd166;
	sample_rom[88][48] = 8'd162;
	sample_rom[88][49] = 8'd156;
	sample_rom[88][50] = 8'd152;
	sample_rom[88][51] = 8'd145;
	sample_rom[88][52] = 8'd143;
	sample_rom[88][53] = 8'd141;
	sample_rom[88][54] = 8'd141;
	sample_rom[88][55] = 8'd142;
	sample_rom[88][56] = 8'd142;
	sample_rom[88][57] = 8'd140;
	sample_rom[88][58] = 8'd139;
	sample_rom[88][59] = 8'd137;
	sample_rom[88][60] = 8'd133;
	sample_rom[88][61] = 8'd129;
	sample_rom[88][62] = 8'd127;
	sample_rom[88][63] = 8'd125;
	sample_rom[89][0] = 8'd131;
	sample_rom[89][1] = 8'd188;
	sample_rom[89][2] = 8'd227;
	sample_rom[89][3] = 8'd247;
	sample_rom[89][4] = 8'd249;
	sample_rom[89][5] = 8'd246;
	sample_rom[89][6] = 8'd243;
	sample_rom[89][7] = 8'd244;
	sample_rom[89][8] = 8'd242;
	sample_rom[89][9] = 8'd240;
	sample_rom[89][10] = 8'd237;
	sample_rom[89][11] = 8'd235;
	sample_rom[89][12] = 8'd233;
	sample_rom[89][13] = 8'd233;
	sample_rom[89][14] = 8'd234;
	sample_rom[89][15] = 8'd235;
	sample_rom[89][16] = 8'd231;
	sample_rom[89][17] = 8'd226;
	sample_rom[89][18] = 8'd223;
	sample_rom[89][19] = 8'd218;
	sample_rom[89][20] = 8'd216;
	sample_rom[89][21] = 8'd217;
	sample_rom[89][22] = 8'd217;
	sample_rom[89][23] = 8'd215;
	sample_rom[89][24] = 8'd209;
	sample_rom[89][25] = 8'd208;
	sample_rom[89][26] = 8'd209;
	sample_rom[89][27] = 8'd203;
	sample_rom[89][28] = 8'd202;
	sample_rom[89][29] = 8'd200;
	sample_rom[89][30] = 8'd198;
	sample_rom[89][31] = 8'd197;
	sample_rom[89][32] = 8'd196;
	sample_rom[89][33] = 8'd199;
	sample_rom[89][34] = 8'd192;
	sample_rom[89][35] = 8'd183;
	sample_rom[89][36] = 8'd182;
	sample_rom[89][37] = 8'd180;
	sample_rom[89][38] = 8'd183;
	sample_rom[89][39] = 8'd177;
	sample_rom[89][40] = 8'd175;
	sample_rom[89][41] = 8'd167;
	sample_rom[89][42] = 8'd164;
	sample_rom[89][43] = 8'd163;
	sample_rom[89][44] = 8'd161;
	sample_rom[89][45] = 8'd165;
	sample_rom[89][46] = 8'd159;
	sample_rom[89][47] = 8'd158;
	sample_rom[89][48] = 8'd156;
	sample_rom[89][49] = 8'd154;
	sample_rom[89][50] = 8'd156;
	sample_rom[89][51] = 8'd148;
	sample_rom[89][52] = 8'd144;
	sample_rom[89][53] = 8'd143;
	sample_rom[89][54] = 8'd143;
	sample_rom[89][55] = 8'd141;
	sample_rom[89][56] = 8'd136;
	sample_rom[89][57] = 8'd132;
	sample_rom[89][58] = 8'd129;
	sample_rom[89][59] = 8'd127;
	sample_rom[89][60] = 8'd127;
	sample_rom[89][61] = 8'd127;
	sample_rom[89][62] = 8'd123;
	sample_rom[89][63] = 8'd126;
	sample_rom[90][0] = 8'd132;
	sample_rom[90][1] = 8'd180;
	sample_rom[90][2] = 8'd217;
	sample_rom[90][3] = 8'd242;
	sample_rom[90][4] = 8'd251;
	sample_rom[90][5] = 8'd253;
	sample_rom[90][6] = 8'd250;
	sample_rom[90][7] = 8'd239;
	sample_rom[90][8] = 8'd224;
	sample_rom[90][9] = 8'd209;
	sample_rom[90][10] = 8'd201;
	sample_rom[90][11] = 8'd194;
	sample_rom[90][12] = 8'd195;
	sample_rom[90][13] = 8'd189;
	sample_rom[90][14] = 8'd187;
	sample_rom[90][15] = 8'd182;
	sample_rom[90][16] = 8'd178;
	sample_rom[90][17] = 8'd170;
	sample_rom[90][18] = 8'd168;
	sample_rom[90][19] = 8'd161;
	sample_rom[90][20] = 8'd158;
	sample_rom[90][21] = 8'd153;
	sample_rom[90][22] = 8'd152;
	sample_rom[90][23] = 8'd153;
	sample_rom[90][24] = 8'd152;
	sample_rom[90][25] = 8'd148;
	sample_rom[90][26] = 8'd135;
	sample_rom[90][27] = 8'd127;
	sample_rom[90][28] = 8'd113;
	sample_rom[90][29] = 8'd105;
	sample_rom[90][30] = 8'd99;
	sample_rom[90][31] = 8'd97;
	sample_rom[90][32] = 8'd100;
	sample_rom[90][33] = 8'd106;
	sample_rom[90][34] = 8'd114;
	sample_rom[90][35] = 8'd122;
	sample_rom[90][36] = 8'd131;
	sample_rom[90][37] = 8'd135;
	sample_rom[90][38] = 8'd141;
	sample_rom[90][39] = 8'd144;
	sample_rom[90][40] = 8'd144;
	sample_rom[90][41] = 8'd142;
	sample_rom[90][42] = 8'd142;
	sample_rom[90][43] = 8'd141;
	sample_rom[90][44] = 8'd145;
	sample_rom[90][45] = 8'd148;
	sample_rom[90][46] = 8'd143;
	sample_rom[90][47] = 8'd134;
	sample_rom[90][48] = 8'd125;
	sample_rom[90][49] = 8'd117;
	sample_rom[90][50] = 8'd111;
	sample_rom[90][51] = 8'd109;
	sample_rom[90][52] = 8'd107;
	sample_rom[90][53] = 8'd104;
	sample_rom[90][54] = 8'd106;
	sample_rom[90][55] = 8'd111;
	sample_rom[90][56] = 8'd118;
	sample_rom[90][57] = 8'd122;
	sample_rom[90][58] = 8'd125;
	sample_rom[90][59] = 8'd128;
	sample_rom[90][60] = 8'd129;
	sample_rom[90][61] = 8'd134;
	sample_rom[90][62] = 8'd136;
	sample_rom[90][63] = 8'd133;
	sample_rom[91][0] = 8'd131;
	sample_rom[91][1] = 8'd178;
	sample_rom[91][2] = 8'd218;
	sample_rom[91][3] = 8'd239;
	sample_rom[91][4] = 8'd247;
	sample_rom[91][5] = 8'd245;
	sample_rom[91][6] = 8'd232;
	sample_rom[91][7] = 8'd216;
	sample_rom[91][8] = 8'd203;
	sample_rom[91][9] = 8'd192;
	sample_rom[91][10] = 8'd186;
	sample_rom[91][11] = 8'd185;
	sample_rom[91][12] = 8'd187;
	sample_rom[91][13] = 8'd190;
	sample_rom[91][14] = 8'd191;
	sample_rom[91][15] = 8'd190;
	sample_rom[91][16] = 8'd182;
	sample_rom[91][17] = 8'd169;
	sample_rom[91][18] = 8'd153;
	sample_rom[91][19] = 8'd131;
	sample_rom[91][20] = 8'd110;
	sample_rom[91][21] = 8'd95;
	sample_rom[91][22] = 8'd87;
	sample_rom[91][23] = 8'd84;
	sample_rom[91][24] = 8'd88;
	sample_rom[91][25] = 8'd94;
	sample_rom[91][26] = 8'd98;
	sample_rom[91][27] = 8'd101;
	sample_rom[91][28] = 8'd101;
	sample_rom[91][29] = 8'd102;
	sample_rom[91][30] = 8'd104;
	sample_rom[91][31] = 8'd104;
	sample_rom[91][32] = 8'd111;
	sample_rom[91][33] = 8'd114;
	sample_rom[91][34] = 8'd121;
	sample_rom[91][35] = 8'd131;
	sample_rom[91][36] = 8'd136;
	sample_rom[91][37] = 8'd145;
	sample_rom[91][38] = 8'd149;
	sample_rom[91][39] = 8'd151;
	sample_rom[91][40] = 8'd148;
	sample_rom[91][41] = 8'd140;
	sample_rom[91][42] = 8'd133;
	sample_rom[91][43] = 8'd121;
	sample_rom[91][44] = 8'd116;
	sample_rom[91][45] = 8'd110;
	sample_rom[91][46] = 8'd108;
	sample_rom[91][47] = 8'd111;
	sample_rom[91][48] = 8'd113;
	sample_rom[91][49] = 8'd111;
	sample_rom[91][50] = 8'd111;
	sample_rom[91][51] = 8'd110;
	sample_rom[91][52] = 8'd111;
	sample_rom[91][53] = 8'd106;
	sample_rom[91][54] = 8'd108;
	sample_rom[91][55] = 8'd109;
	sample_rom[91][56] = 8'd112;
	sample_rom[91][57] = 8'd114;
	sample_rom[91][58] = 8'd111;
	sample_rom[91][59] = 8'd112;
	sample_rom[91][60] = 8'd114;
	sample_rom[91][61] = 8'd117;
	sample_rom[91][62] = 8'd118;
	sample_rom[91][63] = 8'd124;
	sample_rom[92][0] = 8'd132;
	sample_rom[92][1] = 8'd176;
	sample_rom[92][2] = 8'd211;
	sample_rom[92][3] = 8'd232;
	sample_rom[92][4] = 8'd235;
	sample_rom[92][5] = 8'd224;
	sample_rom[92][6] = 8'd201;
	sample_rom[92][7] = 8'd176;
	sample_rom[92][8] = 8'd154;
	sample_rom[92][9] = 8'd139;
	sample_rom[92][10] = 8'd137;
	sample_rom[92][11] = 8'd140;
	sample_rom[92][12] = 8'd153;
	sample_rom[92][13] = 8'd160;
	sample_rom[92][14] = 8'd167;
	sample_rom[92][15] = 8'd171;
	sample_rom[92][16] = 8'd168;
	sample_rom[92][17] = 8'd162;
	sample_rom[92][18] = 8'd156;
	sample_rom[92][19] = 8'd150;
	sample_rom[92][20] = 8'd150;
	sample_rom[92][21] = 8'd153;
	sample_rom[92][22] = 8'd160;
	sample_rom[92][23] = 8'd168;
	sample_rom[92][24] = 8'd176;
	sample_rom[92][25] = 8'd181;
	sample_rom[92][26] = 8'd180;
	sample_rom[92][27] = 8'd173;
	sample_rom[92][28] = 8'd160;
	sample_rom[92][29] = 8'd145;
	sample_rom[92][30] = 8'd130;
	sample_rom[92][31] = 8'd120;
	sample_rom[92][32] = 8'd119;
	sample_rom[92][33] = 8'd123;
	sample_rom[92][34] = 8'd133;
	sample_rom[92][35] = 8'd145;
	sample_rom[92][36] = 8'd154;
	sample_rom[92][37] = 8'd158;
	sample_rom[92][38] = 8'd154;
	sample_rom[92][39] = 8'd145;
	sample_rom[92][40] = 8'd132;
	sample_rom[92][41] = 8'd118;
	sample_rom[92][42] = 8'd106;
	sample_rom[92][43] = 8'd104;
	sample_rom[92][44] = 8'd110;
	sample_rom[92][45] = 8'd121;
	sample_rom[92][46] = 8'd138;
	sample_rom[92][47] = 8'd158;
	sample_rom[92][48] = 8'd174;
	sample_rom[92][49] = 8'd184;
	sample_rom[92][50] = 8'd187;
	sample_rom[92][51] = 8'd184;
	sample_rom[92][52] = 8'd173;
	sample_rom[92][53] = 8'd159;
	sample_rom[92][54] = 8'd140;
	sample_rom[92][55] = 8'd123;
	sample_rom[92][56] = 8'd114;
	sample_rom[92][57] = 8'd108;
	sample_rom[92][58] = 8'd105;
	sample_rom[92][59] = 8'd108;
	sample_rom[92][60] = 8'd113;
	sample_rom[92][61] = 8'd117;
	sample_rom[92][62] = 8'd121;
	sample_rom[92][63] = 8'd126;
	sample_rom[93][0] = 8'd129;
	sample_rom[93][1] = 8'd152;
	sample_rom[93][2] = 8'd170;
	sample_rom[93][3] = 8'd185;
	sample_rom[93][4] = 8'd199;
	sample_rom[93][5] = 8'd207;
	sample_rom[93][6] = 8'd211;
	sample_rom[93][7] = 8'd211;
	sample_rom[93][8] = 8'd208;
	sample_rom[93][9] = 8'd201;
	sample_rom[93][10] = 8'd193;
	sample_rom[93][11] = 8'd181;
	sample_rom[93][12] = 8'd172;
	sample_rom[93][13] = 8'd162;
	sample_rom[93][14] = 8'd155;
	sample_rom[93][15] = 8'd150;
	sample_rom[93][16] = 8'd146;
	sample_rom[93][17] = 8'd143;
	sample_rom[93][18] = 8'd143;
	sample_rom[93][19] = 8'd144;
	sample_rom[93][20] = 8'd144;
	sample_rom[93][21] = 8'd145;
	sample_rom[93][22] = 8'd142;
	sample_rom[93][23] = 8'd143;
	sample_rom[93][24] = 8'd140;
	sample_rom[93][25] = 8'd133;
	sample_rom[93][26] = 8'd130;
	sample_rom[93][27] = 8'd124;
	sample_rom[93][28] = 8'd116;
	sample_rom[93][29] = 8'd110;
	sample_rom[93][30] = 8'd105;
	sample_rom[93][31] = 8'd100;
	sample_rom[93][32] = 8'd99;
	sample_rom[93][33] = 8'd101;
	sample_rom[93][34] = 8'd102;
	sample_rom[93][35] = 8'd107;
	sample_rom[93][36] = 8'd112;
	sample_rom[93][37] = 8'd118;
	sample_rom[93][38] = 8'd126;
	sample_rom[93][39] = 8'd132;
	sample_rom[93][40] = 8'd137;
	sample_rom[93][41] = 8'd140;
	sample_rom[93][42] = 8'd145;
	sample_rom[93][43] = 8'd145;
	sample_rom[93][44] = 8'd146;
	sample_rom[93][45] = 8'd146;
	sample_rom[93][46] = 8'd145;
	sample_rom[93][47] = 8'd146;
	sample_rom[93][48] = 8'd146;
	sample_rom[93][49] = 8'd148;
	sample_rom[93][50] = 8'd152;
	sample_rom[93][51] = 8'd158;
	sample_rom[93][52] = 8'd162;
	sample_rom[93][53] = 8'd171;
	sample_rom[93][54] = 8'd177;
	sample_rom[93][55] = 8'd182;
	sample_rom[93][56] = 8'd187;
	sample_rom[93][57] = 8'd190;
	sample_rom[93][58] = 8'd191;
	sample_rom[93][59] = 8'd186;
	sample_rom[93][60] = 8'd180;
	sample_rom[93][61] = 8'd168;
	sample_rom[93][62] = 8'd157;
	sample_rom[93][63] = 8'd142;
	sample_rom[94][0] = 8'd130;
	sample_rom[94][1] = 8'd137;
	sample_rom[94][2] = 8'd144;
	sample_rom[94][3] = 8'd149;
	sample_rom[94][4] = 8'd156;
	sample_rom[94][5] = 8'd160;
	sample_rom[94][6] = 8'd165;
	sample_rom[94][7] = 8'd169;
	sample_rom[94][8] = 8'd174;
	sample_rom[94][9] = 8'd179;
	sample_rom[94][10] = 8'd185;
	sample_rom[94][11] = 8'd189;
	sample_rom[94][12] = 8'd191;
	sample_rom[94][13] = 8'd195;
	sample_rom[94][14] = 8'd198;
	sample_rom[94][15] = 8'd202;
	sample_rom[94][16] = 8'd204;
	sample_rom[94][17] = 8'd206;
	sample_rom[94][18] = 8'd206;
	sample_rom[94][19] = 8'd208;
	sample_rom[94][20] = 8'd209;
	sample_rom[94][21] = 8'd211;
	sample_rom[94][22] = 8'd211;
	sample_rom[94][23] = 8'd213;
	sample_rom[94][24] = 8'd212;
	sample_rom[94][25] = 8'd213;
	sample_rom[94][26] = 8'd213;
	sample_rom[94][27] = 8'd214;
	sample_rom[94][28] = 8'd214;
	sample_rom[94][29] = 8'd213;
	sample_rom[94][30] = 8'd214;
	sample_rom[94][31] = 8'd213;
	sample_rom[94][32] = 8'd213;
	sample_rom[94][33] = 8'd214;
	sample_rom[94][34] = 8'd213;
	sample_rom[94][35] = 8'd213;
	sample_rom[94][36] = 8'd213;
	sample_rom[94][37] = 8'd212;
	sample_rom[94][38] = 8'd212;
	sample_rom[94][39] = 8'd211;
	sample_rom[94][40] = 8'd212;
	sample_rom[94][41] = 8'd210;
	sample_rom[94][42] = 8'd210;
	sample_rom[94][43] = 8'd208;
	sample_rom[94][44] = 8'd207;
	sample_rom[94][45] = 8'd205;
	sample_rom[94][46] = 8'd205;
	sample_rom[94][47] = 8'd203;
	sample_rom[94][48] = 8'd201;
	sample_rom[94][49] = 8'd198;
	sample_rom[94][50] = 8'd195;
	sample_rom[94][51] = 8'd191;
	sample_rom[94][52] = 8'd188;
	sample_rom[94][53] = 8'd185;
	sample_rom[94][54] = 8'd180;
	sample_rom[94][55] = 8'd174;
	sample_rom[94][56] = 8'd170;
	sample_rom[94][57] = 8'd165;
	sample_rom[94][58] = 8'd160;
	sample_rom[94][59] = 8'd156;
	sample_rom[94][60] = 8'd150;
	sample_rom[94][61] = 8'd145;
	sample_rom[94][62] = 8'd138;
	sample_rom[94][63] = 8'd131;
	sample_rom[95][0] = 8'd132;
	sample_rom[95][1] = 8'd144;
	sample_rom[95][2] = 8'd156;
	sample_rom[95][3] = 8'd164;
	sample_rom[95][4] = 8'd173;
	sample_rom[95][5] = 8'd180;
	sample_rom[95][6] = 8'd187;
	sample_rom[95][7] = 8'd191;
	sample_rom[95][8] = 8'd195;
	sample_rom[95][9] = 8'd199;
	sample_rom[95][10] = 8'd201;
	sample_rom[95][11] = 8'd204;
	sample_rom[95][12] = 8'd205;
	sample_rom[95][13] = 8'd207;
	sample_rom[95][14] = 8'd209;
	sample_rom[95][15] = 8'd212;
	sample_rom[95][16] = 8'd212;
	sample_rom[95][17] = 8'd212;
	sample_rom[95][18] = 8'd212;
	sample_rom[95][19] = 8'd213;
	sample_rom[95][20] = 8'd213;
	sample_rom[95][21] = 8'd213;
	sample_rom[95][22] = 8'd211;
	sample_rom[95][23] = 8'd214;
	sample_rom[95][24] = 8'd212;
	sample_rom[95][25] = 8'd213;
	sample_rom[95][26] = 8'd213;
	sample_rom[95][27] = 8'd214;
	sample_rom[95][28] = 8'd215;
	sample_rom[95][29] = 8'd217;
	sample_rom[95][30] = 8'd218;
	sample_rom[95][31] = 8'd218;
	sample_rom[95][32] = 8'd218;
	sample_rom[95][33] = 8'd217;
	sample_rom[95][34] = 8'd217;
	sample_rom[95][35] = 8'd215;
	sample_rom[95][36] = 8'd215;
	sample_rom[95][37] = 8'd213;
	sample_rom[95][38] = 8'd213;
	sample_rom[95][39] = 8'd211;
	sample_rom[95][40] = 8'd211;
	sample_rom[95][41] = 8'd210;
	sample_rom[95][42] = 8'd211;
	sample_rom[95][43] = 8'd211;
	sample_rom[95][44] = 8'd210;
	sample_rom[95][45] = 8'd210;
	sample_rom[95][46] = 8'd211;
	sample_rom[95][47] = 8'd211;
	sample_rom[95][48] = 8'd210;
	sample_rom[95][49] = 8'd207;
	sample_rom[95][50] = 8'd206;
	sample_rom[95][51] = 8'd204;
	sample_rom[95][52] = 8'd202;
	sample_rom[95][53] = 8'd199;
	sample_rom[95][54] = 8'd197;
	sample_rom[95][55] = 8'd193;
	sample_rom[95][56] = 8'd190;
	sample_rom[95][57] = 8'd186;
	sample_rom[95][58] = 8'd181;
	sample_rom[95][59] = 8'd176;
	sample_rom[95][60] = 8'd167;
	sample_rom[95][61] = 8'd159;
	sample_rom[95][62] = 8'd147;
	sample_rom[95][63] = 8'd138;
	sample_rom[96][0] = 8'd130;
	sample_rom[96][1] = 8'd141;
	sample_rom[96][2] = 8'd152;
	sample_rom[96][3] = 8'd160;
	sample_rom[96][4] = 8'd168;
	sample_rom[96][5] = 8'd174;
	sample_rom[96][6] = 8'd182;
	sample_rom[96][7] = 8'd187;
	sample_rom[96][8] = 8'd192;
	sample_rom[96][9] = 8'd197;
	sample_rom[96][10] = 8'd200;
	sample_rom[96][11] = 8'd202;
	sample_rom[96][12] = 8'd203;
	sample_rom[96][13] = 8'd203;
	sample_rom[96][14] = 8'd204;
	sample_rom[96][15] = 8'd204;
	sample_rom[96][16] = 8'd203;
	sample_rom[96][17] = 8'd203;
	sample_rom[96][18] = 8'd202;
	sample_rom[96][19] = 8'd201;
	sample_rom[96][20] = 8'd201;
	sample_rom[96][21] = 8'd202;
	sample_rom[96][22] = 8'd203;
	sample_rom[96][23] = 8'd204;
	sample_rom[96][24] = 8'd205;
	sample_rom[96][25] = 8'd207;
	sample_rom[96][26] = 8'd207;
	sample_rom[96][27] = 8'd209;
	sample_rom[96][28] = 8'd212;
	sample_rom[96][29] = 8'd212;
	sample_rom[96][30] = 8'd214;
	sample_rom[96][31] = 8'd213;
	sample_rom[96][32] = 8'd214;
	sample_rom[96][33] = 8'd213;
	sample_rom[96][34] = 8'd212;
	sample_rom[96][35] = 8'd212;
	sample_rom[96][36] = 8'd210;
	sample_rom[96][37] = 8'd208;
	sample_rom[96][38] = 8'd207;
	sample_rom[96][39] = 8'd204;
	sample_rom[96][40] = 8'd204;
	sample_rom[96][41] = 8'd202;
	sample_rom[96][42] = 8'd203;
	sample_rom[96][43] = 8'd199;
	sample_rom[96][44] = 8'd200;
	sample_rom[96][45] = 8'd199;
	sample_rom[96][46] = 8'd201;
	sample_rom[96][47] = 8'd201;
	sample_rom[96][48] = 8'd201;
	sample_rom[96][49] = 8'd201;
	sample_rom[96][50] = 8'd201;
	sample_rom[96][51] = 8'd200;
	sample_rom[96][52] = 8'd200;
	sample_rom[96][53] = 8'd198;
	sample_rom[96][54] = 8'd195;
	sample_rom[96][55] = 8'd191;
	sample_rom[96][56] = 8'd188;
	sample_rom[96][57] = 8'd183;
	sample_rom[96][58] = 8'd177;
	sample_rom[96][59] = 8'd171;
	sample_rom[96][60] = 8'd162;
	sample_rom[96][61] = 8'd155;
	sample_rom[96][62] = 8'd144;
	sample_rom[96][63] = 8'd135;
	sample_rom[97][0] = 8'd131;
	sample_rom[97][1] = 8'd154;
	sample_rom[97][2] = 8'd173;
	sample_rom[97][3] = 8'd187;
	sample_rom[97][4] = 8'd193;
	sample_rom[97][5] = 8'd197;
	sample_rom[97][6] = 8'd194;
	sample_rom[97][7] = 8'd193;
	sample_rom[97][8] = 8'd194;
	sample_rom[97][9] = 8'd198;
	sample_rom[97][10] = 8'd201;
	sample_rom[97][11] = 8'd203;
	sample_rom[97][12] = 8'd206;
	sample_rom[97][13] = 8'd206;
	sample_rom[97][14] = 8'd207;
	sample_rom[97][15] = 8'd205;
	sample_rom[97][16] = 8'd206;
	sample_rom[97][17] = 8'd205;
	sample_rom[97][18] = 8'd206;
	sample_rom[97][19] = 8'd208;
	sample_rom[97][20] = 8'd209;
	sample_rom[97][21] = 8'd211;
	sample_rom[97][22] = 8'd210;
	sample_rom[97][23] = 8'd211;
	sample_rom[97][24] = 8'd210;
	sample_rom[97][25] = 8'd211;
	sample_rom[97][26] = 8'd212;
	sample_rom[97][27] = 8'd213;
	sample_rom[97][28] = 8'd214;
	sample_rom[97][29] = 8'd215;
	sample_rom[97][30] = 8'd216;
	sample_rom[97][31] = 8'd216;
	sample_rom[97][32] = 8'd215;
	sample_rom[97][33] = 8'd216;
	sample_rom[97][34] = 8'd215;
	sample_rom[97][35] = 8'd214;
	sample_rom[97][36] = 8'd213;
	sample_rom[97][37] = 8'd211;
	sample_rom[97][38] = 8'd212;
	sample_rom[97][39] = 8'd209;
	sample_rom[97][40] = 8'd210;
	sample_rom[97][41] = 8'd208;
	sample_rom[97][42] = 8'd210;
	sample_rom[97][43] = 8'd209;
	sample_rom[97][44] = 8'd208;
	sample_rom[97][45] = 8'd206;
	sample_rom[97][46] = 8'd205;
	sample_rom[97][47] = 8'd204;
	sample_rom[97][48] = 8'd203;
	sample_rom[97][49] = 8'd203;
	sample_rom[97][50] = 8'd203;
	sample_rom[97][51] = 8'd205;
	sample_rom[97][52] = 8'd203;
	sample_rom[97][53] = 8'd201;
	sample_rom[97][54] = 8'd197;
	sample_rom[97][55] = 8'd193;
	sample_rom[97][56] = 8'd189;
	sample_rom[97][57] = 8'd187;
	sample_rom[97][58] = 8'd191;
	sample_rom[97][59] = 8'd191;
	sample_rom[97][60] = 8'd187;
	sample_rom[97][61] = 8'd180;
	sample_rom[97][62] = 8'd164;
	sample_rom[97][63] = 8'd145;
	sample_rom[98][0] = 8'd132;
	sample_rom[98][1] = 8'd172;
	sample_rom[98][2] = 8'd204;
	sample_rom[98][3] = 8'd218;
	sample_rom[98][4] = 8'd221;
	sample_rom[98][5] = 8'd214;
	sample_rom[98][6] = 8'd205;
	sample_rom[98][7] = 8'd204;
	sample_rom[98][8] = 8'd205;
	sample_rom[98][9] = 8'd204;
	sample_rom[98][10] = 8'd205;
	sample_rom[98][11] = 8'd202;
	sample_rom[98][12] = 8'd201;
	sample_rom[98][13] = 8'd197;
	sample_rom[98][14] = 8'd197;
	sample_rom[98][15] = 8'd198;
	sample_rom[98][16] = 8'd197;
	sample_rom[98][17] = 8'd200;
	sample_rom[98][18] = 8'd205;
	sample_rom[98][19] = 8'd210;
	sample_rom[98][20] = 8'd214;
	sample_rom[98][21] = 8'd223;
	sample_rom[98][22] = 8'd220;
	sample_rom[98][23] = 8'd221;
	sample_rom[98][24] = 8'd218;
	sample_rom[98][25] = 8'd217;
	sample_rom[98][26] = 8'd215;
	sample_rom[98][27] = 8'd214;
	sample_rom[98][28] = 8'd211;
	sample_rom[98][29] = 8'd207;
	sample_rom[98][30] = 8'd201;
	sample_rom[98][31] = 8'd196;
	sample_rom[98][32] = 8'd196;
	sample_rom[98][33] = 8'd201;
	sample_rom[98][34] = 8'd203;
	sample_rom[98][35] = 8'd204;
	sample_rom[98][36] = 8'd208;
	sample_rom[98][37] = 8'd212;
	sample_rom[98][38] = 8'd217;
	sample_rom[98][39] = 8'd219;
	sample_rom[98][40] = 8'd220;
	sample_rom[98][41] = 8'd217;
	sample_rom[98][42] = 8'd219;
	sample_rom[98][43] = 8'd213;
	sample_rom[98][44] = 8'd212;
	sample_rom[98][45] = 8'd207;
	sample_rom[98][46] = 8'd203;
	sample_rom[98][47] = 8'd201;
	sample_rom[98][48] = 8'd194;
	sample_rom[98][49] = 8'd191;
	sample_rom[98][50] = 8'd195;
	sample_rom[98][51] = 8'd199;
	sample_rom[98][52] = 8'd199;
	sample_rom[98][53] = 8'd199;
	sample_rom[98][54] = 8'd194;
	sample_rom[98][55] = 8'd192;
	sample_rom[98][56] = 8'd195;
	sample_rom[98][57] = 8'd205;
	sample_rom[98][58] = 8'd215;
	sample_rom[98][59] = 8'd221;
	sample_rom[98][60] = 8'd216;
	sample_rom[98][61] = 8'd200;
	sample_rom[98][62] = 8'd178;
	sample_rom[98][63] = 8'd153;
	sample_rom[99][0] = 8'd131;
	sample_rom[99][1] = 8'd158;
	sample_rom[99][2] = 8'd179;
	sample_rom[99][3] = 8'd199;
	sample_rom[99][4] = 8'd214;
	sample_rom[99][5] = 8'd225;
	sample_rom[99][6] = 8'd234;
	sample_rom[99][7] = 8'd239;
	sample_rom[99][8] = 8'd243;
	sample_rom[99][9] = 8'd243;
	sample_rom[99][10] = 8'd246;
	sample_rom[99][11] = 8'd246;
	sample_rom[99][12] = 8'd244;
	sample_rom[99][13] = 8'd242;
	sample_rom[99][14] = 8'd240;
	sample_rom[99][15] = 8'd234;
	sample_rom[99][16] = 8'd229;
	sample_rom[99][17] = 8'd218;
	sample_rom[99][18] = 8'd210;
	sample_rom[99][19] = 8'd200;
	sample_rom[99][20] = 8'd192;
	sample_rom[99][21] = 8'd182;
	sample_rom[99][22] = 8'd170;
	sample_rom[99][23] = 8'd166;
	sample_rom[99][24] = 8'd157;
	sample_rom[99][25] = 8'd150;
	sample_rom[99][26] = 8'd146;
	sample_rom[99][27] = 8'd140;
	sample_rom[99][28] = 8'd136;
	sample_rom[99][29] = 8'd133;
	sample_rom[99][30] = 8'd132;
	sample_rom[99][31] = 8'd125;
	sample_rom[99][32] = 8'd123;
	sample_rom[99][33] = 8'd122;
	sample_rom[99][34] = 8'd121;
	sample_rom[99][35] = 8'd121;
	sample_rom[99][36] = 8'd120;
	sample_rom[99][37] = 8'd116;
	sample_rom[99][38] = 8'd118;
	sample_rom[99][39] = 8'd119;
	sample_rom[99][40] = 8'd119;
	sample_rom[99][41] = 8'd122;
	sample_rom[99][42] = 8'd124;
	sample_rom[99][43] = 8'd126;
	sample_rom[99][44] = 8'd132;
	sample_rom[99][45] = 8'd131;
	sample_rom[99][46] = 8'd134;
	sample_rom[99][47] = 8'd135;
	sample_rom[99][48] = 8'd137;
	sample_rom[99][49] = 8'd136;
	sample_rom[99][50] = 8'd137;
	sample_rom[99][51] = 8'd139;
	sample_rom[99][52] = 8'd139;
	sample_rom[99][53] = 8'd140;
	sample_rom[99][54] = 8'd139;
	sample_rom[99][55] = 8'd138;
	sample_rom[99][56] = 8'd139;
	sample_rom[99][57] = 8'd139;
	sample_rom[99][58] = 8'd140;
	sample_rom[99][59] = 8'd135;
	sample_rom[99][60] = 8'd134;
	sample_rom[99][61] = 8'd133;
	sample_rom[99][62] = 8'd129;
	sample_rom[99][63] = 8'd130;
	sample_rom[100][0] = 8'd131;
	sample_rom[100][1] = 8'd175;
	sample_rom[100][2] = 8'd194;
	sample_rom[100][3] = 8'd190;
	sample_rom[100][4] = 8'd186;
	sample_rom[100][5] = 8'd188;
	sample_rom[100][6] = 8'd189;
	sample_rom[100][7] = 8'd186;
	sample_rom[100][8] = 8'd187;
	sample_rom[100][9] = 8'd189;
	sample_rom[100][10] = 8'd194;
	sample_rom[100][11] = 8'd189;
	sample_rom[100][12] = 8'd188;
	sample_rom[100][13] = 8'd188;
	sample_rom[100][14] = 8'd192;
	sample_rom[100][15] = 8'd191;
	sample_rom[100][16] = 8'd189;
	sample_rom[100][17] = 8'd188;
	sample_rom[100][18] = 8'd187;
	sample_rom[100][19] = 8'd187;
	sample_rom[100][20] = 8'd184;
	sample_rom[100][21] = 8'd189;
	sample_rom[100][22] = 8'd191;
	sample_rom[100][23] = 8'd189;
	sample_rom[100][24] = 8'd187;
	sample_rom[100][25] = 8'd186;
	sample_rom[100][26] = 8'd187;
	sample_rom[100][27] = 8'd187;
	sample_rom[100][28] = 8'd187;
	sample_rom[100][29] = 8'd188;
	sample_rom[100][30] = 8'd193;
	sample_rom[100][31] = 8'd191;
	sample_rom[100][32] = 8'd188;
	sample_rom[100][33] = 8'd191;
	sample_rom[100][34] = 8'd191;
	sample_rom[100][35] = 8'd188;
	sample_rom[100][36] = 8'd185;
	sample_rom[100][37] = 8'd185;
	sample_rom[100][38] = 8'd187;
	sample_rom[100][39] = 8'd185;
	sample_rom[100][40] = 8'd186;
	sample_rom[100][41] = 8'd186;
	sample_rom[100][42] = 8'd190;
	sample_rom[100][43] = 8'd187;
	sample_rom[100][44] = 8'd184;
	sample_rom[100][45] = 8'd185;
	sample_rom[100][46] = 8'd188;
	sample_rom[100][47] = 8'd187;
	sample_rom[100][48] = 8'd187;
	sample_rom[100][49] = 8'd188;
	sample_rom[100][50] = 8'd188;
	sample_rom[100][51] = 8'd187;
	sample_rom[100][52] = 8'd187;
	sample_rom[100][53] = 8'd187;
	sample_rom[100][54] = 8'd190;
	sample_rom[100][55] = 8'd187;
	sample_rom[100][56] = 8'd183;
	sample_rom[100][57] = 8'd184;
	sample_rom[100][58] = 8'd187;
	sample_rom[100][59] = 8'd186;
	sample_rom[100][60] = 8'd181;
	sample_rom[100][61] = 8'd183;
	sample_rom[100][62] = 8'd188;
	sample_rom[100][63] = 8'd169;
	sample_rom[101][0] = 8'd131;
	sample_rom[101][1] = 8'd137;
	sample_rom[101][2] = 8'd144;
	sample_rom[101][3] = 8'd149;
	sample_rom[101][4] = 8'd155;
	sample_rom[101][5] = 8'd159;
	sample_rom[101][6] = 8'd164;
	sample_rom[101][7] = 8'd170;
	sample_rom[101][8] = 8'd174;
	sample_rom[101][9] = 8'd180;
	sample_rom[101][10] = 8'd186;
	sample_rom[101][11] = 8'd191;
	sample_rom[101][12] = 8'd196;
	sample_rom[101][13] = 8'd201;
	sample_rom[101][14] = 8'd205;
	sample_rom[101][15] = 8'd210;
	sample_rom[101][16] = 8'd214;
	sample_rom[101][17] = 8'd218;
	sample_rom[101][18] = 8'd220;
	sample_rom[101][19] = 8'd223;
	sample_rom[101][20] = 8'd226;
	sample_rom[101][21] = 8'd230;
	sample_rom[101][22] = 8'd232;
	sample_rom[101][23] = 8'd235;
	sample_rom[101][24] = 8'd236;
	sample_rom[101][25] = 8'd239;
	sample_rom[101][26] = 8'd240;
	sample_rom[101][27] = 8'd242;
	sample_rom[101][28] = 8'd243;
	sample_rom[101][29] = 8'd244;
	sample_rom[101][30] = 8'd245;
	sample_rom[101][31] = 8'd245;
	sample_rom[101][32] = 8'd245;
	sample_rom[101][33] = 8'd245;
	sample_rom[101][34] = 8'd244;
	sample_rom[101][35] = 8'd243;
	sample_rom[101][36] = 8'd242;
	sample_rom[101][37] = 8'd240;
	sample_rom[101][38] = 8'd239;
	sample_rom[101][39] = 8'd236;
	sample_rom[101][40] = 8'd235;
	sample_rom[101][41] = 8'd232;
	sample_rom[101][42] = 8'd230;
	sample_rom[101][43] = 8'd226;
	sample_rom[101][44] = 8'd223;
	sample_rom[101][45] = 8'd220;
	sample_rom[101][46] = 8'd218;
	sample_rom[101][47] = 8'd214;
	sample_rom[101][48] = 8'd210;
	sample_rom[101][49] = 8'd205;
	sample_rom[101][50] = 8'd201;
	sample_rom[101][51] = 8'd196;
	sample_rom[101][52] = 8'd191;
	sample_rom[101][53] = 8'd186;
	sample_rom[101][54] = 8'd180;
	sample_rom[101][55] = 8'd174;
	sample_rom[101][56] = 8'd170;
	sample_rom[101][57] = 8'd164;
	sample_rom[101][58] = 8'd159;
	sample_rom[101][59] = 8'd155;
	sample_rom[101][60] = 8'd149;
	sample_rom[101][61] = 8'd144;
	sample_rom[101][62] = 8'd137;
	sample_rom[101][63] = 8'd131;
	sample_rom[102][0] = 8'd130;
	sample_rom[102][1] = 8'd163;
	sample_rom[102][2] = 8'd191;
	sample_rom[102][3] = 8'd213;
	sample_rom[102][4] = 8'd230;
	sample_rom[102][5] = 8'd239;
	sample_rom[102][6] = 8'd243;
	sample_rom[102][7] = 8'd241;
	sample_rom[102][8] = 8'd233;
	sample_rom[102][9] = 8'd223;
	sample_rom[102][10] = 8'd206;
	sample_rom[102][11] = 8'd189;
	sample_rom[102][12] = 8'd167;
	sample_rom[102][13] = 8'd146;
	sample_rom[102][14] = 8'd126;
	sample_rom[102][15] = 8'd110;
	sample_rom[102][16] = 8'd95;
	sample_rom[102][17] = 8'd84;
	sample_rom[102][18] = 8'd81;
	sample_rom[102][19] = 8'd78;
	sample_rom[102][20] = 8'd79;
	sample_rom[102][21] = 8'd83;
	sample_rom[102][22] = 8'd90;
	sample_rom[102][23] = 8'd96;
	sample_rom[102][24] = 8'd101;
	sample_rom[102][25] = 8'd113;
	sample_rom[102][26] = 8'd119;
	sample_rom[102][27] = 8'd126;
	sample_rom[102][28] = 8'd130;
	sample_rom[102][29] = 8'd133;
	sample_rom[102][30] = 8'd130;
	sample_rom[102][31] = 8'd129;
	sample_rom[102][32] = 8'd125;
	sample_rom[102][33] = 8'd122;
	sample_rom[102][34] = 8'd118;
	sample_rom[102][35] = 8'd114;
	sample_rom[102][36] = 8'd112;
	sample_rom[102][37] = 8'd110;
	sample_rom[102][38] = 8'd108;
	sample_rom[102][39] = 8'd110;
	sample_rom[102][40] = 8'd113;
	sample_rom[102][41] = 8'd120;
	sample_rom[102][42] = 8'd127;
	sample_rom[102][43] = 8'd133;
	sample_rom[102][44] = 8'd141;
	sample_rom[102][45] = 8'd149;
	sample_rom[102][46] = 8'd155;
	sample_rom[102][47] = 8'd158;
	sample_rom[102][48] = 8'd160;
	sample_rom[102][49] = 8'd160;
	sample_rom[102][50] = 8'd159;
	sample_rom[102][51] = 8'd158;
	sample_rom[102][52] = 8'd154;
	sample_rom[102][53] = 8'd147;
	sample_rom[102][54] = 8'd139;
	sample_rom[102][55] = 8'd133;
	sample_rom[102][56] = 8'd127;
	sample_rom[102][57] = 8'd123;
	sample_rom[102][58] = 8'd121;
	sample_rom[102][59] = 8'd123;
	sample_rom[102][60] = 8'd125;
	sample_rom[102][61] = 8'd126;
	sample_rom[102][62] = 8'd126;
	sample_rom[102][63] = 8'd129;
	sample_rom[103][0] = 8'd128;
	sample_rom[103][1] = 8'd208;
	sample_rom[103][2] = 8'd235;
	sample_rom[103][3] = 8'd232;
	sample_rom[103][4] = 8'd217;
	sample_rom[103][5] = 8'd220;
	sample_rom[103][6] = 8'd229;
	sample_rom[103][7] = 8'd231;
	sample_rom[103][8] = 8'd212;
	sample_rom[103][9] = 8'd176;
	sample_rom[103][10] = 8'd137;
	sample_rom[103][11] = 8'd120;
	sample_rom[103][12] = 8'd123;
	sample_rom[103][13] = 8'd130;
	sample_rom[103][14] = 8'd128;
	sample_rom[103][15] = 8'd125;
	sample_rom[103][16] = 8'd125;
	sample_rom[103][17] = 8'd130;
	sample_rom[103][18] = 8'd133;
	sample_rom[103][19] = 8'd128;
	sample_rom[103][20] = 8'd125;
	sample_rom[103][21] = 8'd130;
	sample_rom[103][22] = 8'd129;
	sample_rom[103][23] = 8'd128;
	sample_rom[103][24] = 8'd129;
	sample_rom[103][25] = 8'd130;
	sample_rom[103][26] = 8'd131;
	sample_rom[103][27] = 8'd129;
	sample_rom[103][28] = 8'd128;
	sample_rom[103][29] = 8'd130;
	sample_rom[103][30] = 8'd130;
	sample_rom[103][31] = 8'd128;
	sample_rom[103][32] = 8'd126;
	sample_rom[103][33] = 8'd130;
	sample_rom[103][34] = 8'd129;
	sample_rom[103][35] = 8'd127;
	sample_rom[103][36] = 8'd129;
	sample_rom[103][37] = 8'd129;
	sample_rom[103][38] = 8'd131;
	sample_rom[103][39] = 8'd127;
	sample_rom[103][40] = 8'd129;
	sample_rom[103][41] = 8'd134;
	sample_rom[103][42] = 8'd131;
	sample_rom[103][43] = 8'd127;
	sample_rom[103][44] = 8'd125;
	sample_rom[103][45] = 8'd130;
	sample_rom[103][46] = 8'd129;
	sample_rom[103][47] = 8'd127;
	sample_rom[103][48] = 8'd128;
	sample_rom[103][49] = 8'd131;
	sample_rom[103][50] = 8'd133;
	sample_rom[103][51] = 8'd131;
	sample_rom[103][52] = 8'd128;
	sample_rom[103][53] = 8'd129;
	sample_rom[103][54] = 8'd132;
	sample_rom[103][55] = 8'd128;
	sample_rom[103][56] = 8'd130;
	sample_rom[103][57] = 8'd127;
	sample_rom[103][58] = 8'd126;
	sample_rom[103][59] = 8'd126;
	sample_rom[103][60] = 8'd126;
	sample_rom[103][61] = 8'd125;
	sample_rom[103][62] = 8'd132;
	sample_rom[103][63] = 8'd128;
	sample_rom[104][0] = 8'd132;
	sample_rom[104][1] = 8'd219;
	sample_rom[104][2] = 8'd250;
	sample_rom[104][3] = 8'd240;
	sample_rom[104][4] = 8'd233;
	sample_rom[104][5] = 8'd241;
	sample_rom[104][6] = 8'd239;
	sample_rom[104][7] = 8'd231;
	sample_rom[104][8] = 8'd228;
	sample_rom[104][9] = 8'd233;
	sample_rom[104][10] = 8'd239;
	sample_rom[104][11] = 8'd233;
	sample_rom[104][12] = 8'd227;
	sample_rom[104][13] = 8'd226;
	sample_rom[104][14] = 8'd225;
	sample_rom[104][15] = 8'd221;
	sample_rom[104][16] = 8'd217;
	sample_rom[104][17] = 8'd219;
	sample_rom[104][18] = 8'd214;
	sample_rom[104][19] = 8'd211;
	sample_rom[104][20] = 8'd205;
	sample_rom[104][21] = 8'd207;
	sample_rom[104][22] = 8'd206;
	sample_rom[104][23] = 8'd206;
	sample_rom[104][24] = 8'd205;
	sample_rom[104][25] = 8'd204;
	sample_rom[104][26] = 8'd200;
	sample_rom[104][27] = 8'd194;
	sample_rom[104][28] = 8'd191;
	sample_rom[104][29] = 8'd192;
	sample_rom[104][30] = 8'd197;
	sample_rom[104][31] = 8'd192;
	sample_rom[104][32] = 8'd189;
	sample_rom[104][33] = 8'd189;
	sample_rom[104][34] = 8'd186;
	sample_rom[104][35] = 8'd179;
	sample_rom[104][36] = 8'd181;
	sample_rom[104][37] = 8'd175;
	sample_rom[104][38] = 8'd177;
	sample_rom[104][39] = 8'd172;
	sample_rom[104][40] = 8'd168;
	sample_rom[104][41] = 8'd169;
	sample_rom[104][42] = 8'd170;
	sample_rom[104][43] = 8'd165;
	sample_rom[104][44] = 8'd166;
	sample_rom[104][45] = 8'd163;
	sample_rom[104][46] = 8'd164;
	sample_rom[104][47] = 8'd156;
	sample_rom[104][48] = 8'd156;
	sample_rom[104][49] = 8'd156;
	sample_rom[104][50] = 8'd153;
	sample_rom[104][51] = 8'd151;
	sample_rom[104][52] = 8'd151;
	sample_rom[104][53] = 8'd149;
	sample_rom[104][54] = 8'd143;
	sample_rom[104][55] = 8'd141;
	sample_rom[104][56] = 8'd139;
	sample_rom[104][57] = 8'd140;
	sample_rom[104][58] = 8'd141;
	sample_rom[104][59] = 8'd141;
	sample_rom[104][60] = 8'd137;
	sample_rom[104][61] = 8'd136;
	sample_rom[104][62] = 8'd133;
	sample_rom[104][63] = 8'd129;
	sample_rom[105][0] = 8'd130;
	sample_rom[105][1] = 8'd176;
	sample_rom[105][2] = 8'd206;
	sample_rom[105][3] = 8'd219;
	sample_rom[105][4] = 8'd216;
	sample_rom[105][5] = 8'd206;
	sample_rom[105][6] = 8'd199;
	sample_rom[105][7] = 8'd198;
	sample_rom[105][8] = 8'd208;
	sample_rom[105][9] = 8'd222;
	sample_rom[105][10] = 8'd230;
	sample_rom[105][11] = 8'd235;
	sample_rom[105][12] = 8'd230;
	sample_rom[105][13] = 8'd225;
	sample_rom[105][14] = 8'd218;
	sample_rom[105][15] = 8'd209;
	sample_rom[105][16] = 8'd208;
	sample_rom[105][17] = 8'd202;
	sample_rom[105][18] = 8'd200;
	sample_rom[105][19] = 8'd191;
	sample_rom[105][20] = 8'd185;
	sample_rom[105][21] = 8'd176;
	sample_rom[105][22] = 8'd166;
	sample_rom[105][23] = 8'd160;
	sample_rom[105][24] = 8'd156;
	sample_rom[105][25] = 8'd148;
	sample_rom[105][26] = 8'd143;
	sample_rom[105][27] = 8'd140;
	sample_rom[105][28] = 8'd135;
	sample_rom[105][29] = 8'd135;
	sample_rom[105][30] = 8'd134;
	sample_rom[105][31] = 8'd130;
	sample_rom[105][32] = 8'd126;
	sample_rom[105][33] = 8'd123;
	sample_rom[105][34] = 8'd119;
	sample_rom[105][35] = 8'd120;
	sample_rom[105][36] = 8'd122;
	sample_rom[105][37] = 8'd120;
	sample_rom[105][38] = 8'd121;
	sample_rom[105][39] = 8'd117;
	sample_rom[105][40] = 8'd117;
	sample_rom[105][41] = 8'd115;
	sample_rom[105][42] = 8'd118;
	sample_rom[105][43] = 8'd121;
	sample_rom[105][44] = 8'd125;
	sample_rom[105][45] = 8'd128;
	sample_rom[105][46] = 8'd129;
	sample_rom[105][47] = 8'd131;
	sample_rom[105][48] = 8'd132;
	sample_rom[105][49] = 8'd130;
	sample_rom[105][50] = 8'd133;
	sample_rom[105][51] = 8'd132;
	sample_rom[105][52] = 8'd138;
	sample_rom[105][53] = 8'd138;
	sample_rom[105][54] = 8'd140;
	sample_rom[105][55] = 8'd136;
	sample_rom[105][56] = 8'd136;
	sample_rom[105][57] = 8'd135;
	sample_rom[105][58] = 8'd136;
	sample_rom[105][59] = 8'd135;
	sample_rom[105][60] = 8'd133;
	sample_rom[105][61] = 8'd133;
	sample_rom[105][62] = 8'd128;
	sample_rom[105][63] = 8'd132;
	sample_rom[106][0] = 8'd130;
	sample_rom[106][1] = 8'd141;
	sample_rom[106][2] = 8'd150;
	sample_rom[106][3] = 8'd154;
	sample_rom[106][4] = 8'd157;
	sample_rom[106][5] = 8'd155;
	sample_rom[106][6] = 8'd154;
	sample_rom[106][7] = 8'd154;
	sample_rom[106][8] = 8'd156;
	sample_rom[106][9] = 8'd162;
	sample_rom[106][10] = 8'd172;
	sample_rom[106][11] = 8'd181;
	sample_rom[106][12] = 8'd189;
	sample_rom[106][13] = 8'd195;
	sample_rom[106][14] = 8'd199;
	sample_rom[106][15] = 8'd199;
	sample_rom[106][16] = 8'd197;
	sample_rom[106][17] = 8'd194;
	sample_rom[106][18] = 8'd193;
	sample_rom[106][19] = 8'd196;
	sample_rom[106][20] = 8'd200;
	sample_rom[106][21] = 8'd209;
	sample_rom[106][22] = 8'd216;
	sample_rom[106][23] = 8'd223;
	sample_rom[106][24] = 8'd225;
	sample_rom[106][25] = 8'd225;
	sample_rom[106][26] = 8'd222;
	sample_rom[106][27] = 8'd219;
	sample_rom[106][28] = 8'd215;
	sample_rom[106][29] = 8'd213;
	sample_rom[106][30] = 8'd214;
	sample_rom[106][31] = 8'd218;
	sample_rom[106][32] = 8'd223;
	sample_rom[106][33] = 8'd228;
	sample_rom[106][34] = 8'd230;
	sample_rom[106][35] = 8'd230;
	sample_rom[106][36] = 8'd227;
	sample_rom[106][37] = 8'd221;
	sample_rom[106][38] = 8'd214;
	sample_rom[106][39] = 8'd208;
	sample_rom[106][40] = 8'd205;
	sample_rom[106][41] = 8'd204;
	sample_rom[106][42] = 8'd208;
	sample_rom[106][43] = 8'd209;
	sample_rom[106][44] = 8'd212;
	sample_rom[106][45] = 8'd211;
	sample_rom[106][46] = 8'd209;
	sample_rom[106][47] = 8'd202;
	sample_rom[106][48] = 8'd194;
	sample_rom[106][49] = 8'd184;
	sample_rom[106][50] = 8'd177;
	sample_rom[106][51] = 8'd173;
	sample_rom[106][52] = 8'd172;
	sample_rom[106][53] = 8'd173;
	sample_rom[106][54] = 8'd174;
	sample_rom[106][55] = 8'd173;
	sample_rom[106][56] = 8'd171;
	sample_rom[106][57] = 8'd165;
	sample_rom[106][58] = 8'd156;
	sample_rom[106][59] = 8'd148;
	sample_rom[106][60] = 8'd138;
	sample_rom[106][61] = 8'd132;
	sample_rom[106][62] = 8'd126;
	sample_rom[106][63] = 8'd125;
	sample_rom[107][0] = 8'd130;
	sample_rom[107][1] = 8'd144;
	sample_rom[107][2] = 8'd154;
	sample_rom[107][3] = 8'd160;
	sample_rom[107][4] = 8'd162;
	sample_rom[107][5] = 8'd163;
	sample_rom[107][6] = 8'd164;
	sample_rom[107][7] = 8'd167;
	sample_rom[107][8] = 8'd172;
	sample_rom[107][9] = 8'd181;
	sample_rom[107][10] = 8'd192;
	sample_rom[107][11] = 8'd203;
	sample_rom[107][12] = 8'd209;
	sample_rom[107][13] = 8'd212;
	sample_rom[107][14] = 8'd210;
	sample_rom[107][15] = 8'd207;
	sample_rom[107][16] = 8'd203;
	sample_rom[107][17] = 8'd202;
	sample_rom[107][18] = 8'd204;
	sample_rom[107][19] = 8'd208;
	sample_rom[107][20] = 8'd213;
	sample_rom[107][21] = 8'd218;
	sample_rom[107][22] = 8'd219;
	sample_rom[107][23] = 8'd216;
	sample_rom[107][24] = 8'd209;
	sample_rom[107][25] = 8'd201;
	sample_rom[107][26] = 8'd192;
	sample_rom[107][27] = 8'd185;
	sample_rom[107][28] = 8'd183;
	sample_rom[107][29] = 8'd185;
	sample_rom[107][30] = 8'd187;
	sample_rom[107][31] = 8'd187;
	sample_rom[107][32] = 8'd184;
	sample_rom[107][33] = 8'd177;
	sample_rom[107][34] = 8'd167;
	sample_rom[107][35] = 8'd157;
	sample_rom[107][36] = 8'd148;
	sample_rom[107][37] = 8'd140;
	sample_rom[107][38] = 8'd139;
	sample_rom[107][39] = 8'd139;
	sample_rom[107][40] = 8'd141;
	sample_rom[107][41] = 8'd142;
	sample_rom[107][42] = 8'd140;
	sample_rom[107][43] = 8'd132;
	sample_rom[107][44] = 8'd124;
	sample_rom[107][45] = 8'd116;
	sample_rom[107][46] = 8'd109;
	sample_rom[107][47] = 8'd106;
	sample_rom[107][48] = 8'd107;
	sample_rom[107][49] = 8'd111;
	sample_rom[107][50] = 8'd116;
	sample_rom[107][51] = 8'd119;
	sample_rom[107][52] = 8'd119;
	sample_rom[107][53] = 8'd116;
	sample_rom[107][54] = 8'd111;
	sample_rom[107][55] = 8'd106;
	sample_rom[107][56] = 8'd102;
	sample_rom[107][57] = 8'd104;
	sample_rom[107][58] = 8'd109;
	sample_rom[107][59] = 8'd118;
	sample_rom[107][60] = 8'd126;
	sample_rom[107][61] = 8'd131;
	sample_rom[107][62] = 8'd132;
	sample_rom[107][63] = 8'd131;
	sample_rom[108][0] = 8'd130;
	sample_rom[108][1] = 8'd147;
	sample_rom[108][2] = 8'd159;
	sample_rom[108][3] = 8'd165;
	sample_rom[108][4] = 8'd168;
	sample_rom[108][5] = 8'd172;
	sample_rom[108][6] = 8'd174;
	sample_rom[108][7] = 8'd180;
	sample_rom[108][8] = 8'd190;
	sample_rom[108][9] = 8'd201;
	sample_rom[108][10] = 8'd213;
	sample_rom[108][11] = 8'd221;
	sample_rom[108][12] = 8'd224;
	sample_rom[108][13] = 8'd223;
	sample_rom[108][14] = 8'd220;
	sample_rom[108][15] = 8'd216;
	sample_rom[108][16] = 8'd213;
	sample_rom[108][17] = 8'd215;
	sample_rom[108][18] = 8'd219;
	sample_rom[108][19] = 8'd223;
	sample_rom[108][20] = 8'd223;
	sample_rom[108][21] = 8'd220;
	sample_rom[108][22] = 8'd210;
	sample_rom[108][23] = 8'd199;
	sample_rom[108][24] = 8'd187;
	sample_rom[108][25] = 8'd176;
	sample_rom[108][26] = 8'd171;
	sample_rom[108][27] = 8'd168;
	sample_rom[108][28] = 8'd165;
	sample_rom[108][29] = 8'd161;
	sample_rom[108][30] = 8'd154;
	sample_rom[108][31] = 8'd141;
	sample_rom[108][32] = 8'd126;
	sample_rom[108][33] = 8'd110;
	sample_rom[108][34] = 8'd97;
	sample_rom[108][35] = 8'd91;
	sample_rom[108][36] = 8'd88;
	sample_rom[108][37] = 8'd84;
	sample_rom[108][38] = 8'd82;
	sample_rom[108][39] = 8'd76;
	sample_rom[108][40] = 8'd66;
	sample_rom[108][41] = 8'd55;
	sample_rom[108][42] = 8'd43;
	sample_rom[108][43] = 8'd35;
	sample_rom[108][44] = 8'd32;
	sample_rom[108][45] = 8'd34;
	sample_rom[108][46] = 8'd36;
	sample_rom[108][47] = 8'd41;
	sample_rom[108][48] = 8'd43;
	sample_rom[108][49] = 8'd41;
	sample_rom[108][50] = 8'd37;
	sample_rom[108][51] = 8'd34;
	sample_rom[108][52] = 8'd34;
	sample_rom[108][53] = 8'd36;
	sample_rom[108][54] = 8'd46;
	sample_rom[108][55] = 8'd57;
	sample_rom[108][56] = 8'd69;
	sample_rom[108][57] = 8'd80;
	sample_rom[108][58] = 8'd85;
	sample_rom[108][59] = 8'd89;
	sample_rom[108][60] = 8'd91;
	sample_rom[108][61] = 8'd95;
	sample_rom[108][62] = 8'd102;
	sample_rom[108][63] = 8'd115;
	sample_rom[109][0] = 8'd130;
	sample_rom[109][1] = 8'd150;
	sample_rom[109][2] = 8'd163;
	sample_rom[109][3] = 8'd171;
	sample_rom[109][4] = 8'd176;
	sample_rom[109][5] = 8'd180;
	sample_rom[109][6] = 8'd184;
	sample_rom[109][7] = 8'd192;
	sample_rom[109][8] = 8'd204;
	sample_rom[109][9] = 8'd215;
	sample_rom[109][10] = 8'd223;
	sample_rom[109][11] = 8'd226;
	sample_rom[109][12] = 8'd223;
	sample_rom[109][13] = 8'd216;
	sample_rom[109][14] = 8'd209;
	sample_rom[109][15] = 8'd203;
	sample_rom[109][16] = 8'd202;
	sample_rom[109][17] = 8'd203;
	sample_rom[109][18] = 8'd201;
	sample_rom[109][19] = 8'd198;
	sample_rom[109][20] = 8'd188;
	sample_rom[109][21] = 8'd172;
	sample_rom[109][22] = 8'd156;
	sample_rom[109][23] = 8'd144;
	sample_rom[109][24] = 8'd134;
	sample_rom[109][25] = 8'd128;
	sample_rom[109][26] = 8'd125;
	sample_rom[109][27] = 8'd121;
	sample_rom[109][28] = 8'd114;
	sample_rom[109][29] = 8'd103;
	sample_rom[109][30] = 8'd91;
	sample_rom[109][31] = 8'd78;
	sample_rom[109][32] = 8'd70;
	sample_rom[109][33] = 8'd69;
	sample_rom[109][34] = 8'd71;
	sample_rom[109][35] = 8'd77;
	sample_rom[109][36] = 8'd80;
	sample_rom[109][37] = 8'd78;
	sample_rom[109][38] = 8'd74;
	sample_rom[109][39] = 8'd69;
	sample_rom[109][40] = 8'd68;
	sample_rom[109][41] = 8'd72;
	sample_rom[109][42] = 8'd81;
	sample_rom[109][43] = 8'd93;
	sample_rom[109][44] = 8'd102;
	sample_rom[109][45] = 8'd108;
	sample_rom[109][46] = 8'd111;
	sample_rom[109][47] = 8'd109;
	sample_rom[109][48] = 8'd108;
	sample_rom[109][49] = 8'd109;
	sample_rom[109][50] = 8'd117;
	sample_rom[109][51] = 8'd127;
	sample_rom[109][52] = 8'd137;
	sample_rom[109][53] = 8'd143;
	sample_rom[109][54] = 8'd145;
	sample_rom[109][55] = 8'd141;
	sample_rom[109][56] = 8'd134;
	sample_rom[109][57] = 8'd129;
	sample_rom[109][58] = 8'd130;
	sample_rom[109][59] = 8'd134;
	sample_rom[109][60] = 8'd139;
	sample_rom[109][61] = 8'd143;
	sample_rom[109][62] = 8'd142;
	sample_rom[109][63] = 8'd136;
	sample_rom[110][0] = 8'd130;
	sample_rom[110][1] = 8'd152;
	sample_rom[110][2] = 8'd167;
	sample_rom[110][3] = 8'd177;
	sample_rom[110][4] = 8'd182;
	sample_rom[110][5] = 8'd187;
	sample_rom[110][6] = 8'd192;
	sample_rom[110][7] = 8'd204;
	sample_rom[110][8] = 8'd216;
	sample_rom[110][9] = 8'd227;
	sample_rom[110][10] = 8'd232;
	sample_rom[110][11] = 8'd229;
	sample_rom[110][12] = 8'd221;
	sample_rom[110][13] = 8'd209;
	sample_rom[110][14] = 8'd201;
	sample_rom[110][15] = 8'd195;
	sample_rom[110][16] = 8'd194;
	sample_rom[110][17] = 8'd189;
	sample_rom[110][18] = 8'd180;
	sample_rom[110][19] = 8'd164;
	sample_rom[110][20] = 8'd145;
	sample_rom[110][21] = 8'd123;
	sample_rom[110][22] = 8'd106;
	sample_rom[110][23] = 8'd97;
	sample_rom[110][24] = 8'd91;
	sample_rom[110][25] = 8'd84;
	sample_rom[110][26] = 8'd76;
	sample_rom[110][27] = 8'd63;
	sample_rom[110][28] = 8'd49;
	sample_rom[110][29] = 8'd35;
	sample_rom[110][30] = 8'd28;
	sample_rom[110][31] = 8'd28;
	sample_rom[110][32] = 8'd34;
	sample_rom[110][33] = 8'd41;
	sample_rom[110][34] = 8'd48;
	sample_rom[110][35] = 8'd51;
	sample_rom[110][36] = 8'd51;
	sample_rom[110][37] = 8'd52;
	sample_rom[110][38] = 8'd60;
	sample_rom[110][39] = 8'd74;
	sample_rom[110][40] = 8'd95;
	sample_rom[110][41] = 8'd113;
	sample_rom[110][42] = 8'd131;
	sample_rom[110][43] = 8'd142;
	sample_rom[110][44] = 8'd150;
	sample_rom[110][45] = 8'd155;
	sample_rom[110][46] = 8'd165;
	sample_rom[110][47] = 8'd179;
	sample_rom[110][48] = 8'd197;
	sample_rom[110][49] = 8'd212;
	sample_rom[110][50] = 8'd222;
	sample_rom[110][51] = 8'd224;
	sample_rom[110][52] = 8'd222;
	sample_rom[110][53] = 8'd216;
	sample_rom[110][54] = 8'd212;
	sample_rom[110][55] = 8'd212;
	sample_rom[110][56] = 8'd215;
	sample_rom[110][57] = 8'd214;
	sample_rom[110][58] = 8'd210;
	sample_rom[110][59] = 8'd197;
	sample_rom[110][60] = 8'd179;
	sample_rom[110][61] = 8'd159;
	sample_rom[110][62] = 8'd143;
	sample_rom[110][63] = 8'd134;
	sample_rom[111][0] = 8'd130;
	sample_rom[111][1] = 8'd155;
	sample_rom[111][2] = 8'd171;
	sample_rom[111][3] = 8'd182;
	sample_rom[111][4] = 8'd188;
	sample_rom[111][5] = 8'd193;
	sample_rom[111][6] = 8'd201;
	sample_rom[111][7] = 8'd212;
	sample_rom[111][8] = 8'd223;
	sample_rom[111][9] = 8'd229;
	sample_rom[111][10] = 8'd226;
	sample_rom[111][11] = 8'd216;
	sample_rom[111][12] = 8'd202;
	sample_rom[111][13] = 8'd188;
	sample_rom[111][14] = 8'd179;
	sample_rom[111][15] = 8'd174;
	sample_rom[111][16] = 8'd167;
	sample_rom[111][17] = 8'd155;
	sample_rom[111][18] = 8'd136;
	sample_rom[111][19] = 8'd113;
	sample_rom[111][20] = 8'd95;
	sample_rom[111][21] = 8'd81;
	sample_rom[111][22] = 8'd74;
	sample_rom[111][23] = 8'd73;
	sample_rom[111][24] = 8'd71;
	sample_rom[111][25] = 8'd65;
	sample_rom[111][26] = 8'd56;
	sample_rom[111][27] = 8'd49;
	sample_rom[111][28] = 8'd46;
	sample_rom[111][29] = 8'd52;
	sample_rom[111][30] = 8'd65;
	sample_rom[111][31] = 8'd79;
	sample_rom[111][32] = 8'd92;
	sample_rom[111][33] = 8'd98;
	sample_rom[111][34] = 8'd100;
	sample_rom[111][35] = 8'd105;
	sample_rom[111][36] = 8'd115;
	sample_rom[111][37] = 8'd128;
	sample_rom[111][38] = 8'd146;
	sample_rom[111][39] = 8'd160;
	sample_rom[111][40] = 8'd167;
	sample_rom[111][41] = 8'd166;
	sample_rom[111][42] = 8'd162;
	sample_rom[111][43] = 8'd161;
	sample_rom[111][44] = 8'd164;
	sample_rom[111][45] = 8'd169;
	sample_rom[111][46] = 8'd174;
	sample_rom[111][47] = 8'd176;
	sample_rom[111][48] = 8'd168;
	sample_rom[111][49] = 8'd155;
	sample_rom[111][50] = 8'd145;
	sample_rom[111][51] = 8'd137;
	sample_rom[111][52] = 8'd135;
	sample_rom[111][53] = 8'd139;
	sample_rom[111][54] = 8'd140;
	sample_rom[111][55] = 8'd136;
	sample_rom[111][56] = 8'd127;
	sample_rom[111][57] = 8'd117;
	sample_rom[111][58] = 8'd112;
	sample_rom[111][59] = 8'd113;
	sample_rom[111][60] = 8'd118;
	sample_rom[111][61] = 8'd127;
	sample_rom[111][62] = 8'd134;
	sample_rom[111][63] = 8'd132;
	sample_rom[112][0] = 8'd130;
	sample_rom[112][1] = 8'd158;
	sample_rom[112][2] = 8'd174;
	sample_rom[112][3] = 8'd186;
	sample_rom[112][4] = 8'd193;
	sample_rom[112][5] = 8'd198;
	sample_rom[112][6] = 8'd208;
	sample_rom[112][7] = 8'd221;
	sample_rom[112][8] = 8'd229;
	sample_rom[112][9] = 8'd230;
	sample_rom[112][10] = 8'd220;
	sample_rom[112][11] = 8'd202;
	sample_rom[112][12] = 8'd185;
	sample_rom[112][13] = 8'd171;
	sample_rom[112][14] = 8'd160;
	sample_rom[112][15] = 8'd151;
	sample_rom[112][16] = 8'd136;
	sample_rom[112][17] = 8'd112;
	sample_rom[112][18] = 8'd89;
	sample_rom[112][19] = 8'd65;
	sample_rom[112][20] = 8'd50;
	sample_rom[112][21] = 8'd47;
	sample_rom[112][22] = 8'd46;
	sample_rom[112][23] = 8'd44;
	sample_rom[112][24] = 8'd40;
	sample_rom[112][25] = 8'd34;
	sample_rom[112][26] = 8'd34;
	sample_rom[112][27] = 8'd42;
	sample_rom[112][28] = 8'd59;
	sample_rom[112][29] = 8'd82;
	sample_rom[112][30] = 8'd103;
	sample_rom[112][31] = 8'd118;
	sample_rom[112][32] = 8'd130;
	sample_rom[112][33] = 8'd143;
	sample_rom[112][34] = 8'd157;
	sample_rom[112][35] = 8'd178;
	sample_rom[112][36] = 8'd201;
	sample_rom[112][37] = 8'd216;
	sample_rom[112][38] = 8'd223;
	sample_rom[112][39] = 8'd223;
	sample_rom[112][40] = 8'd216;
	sample_rom[112][41] = 8'd211;
	sample_rom[112][42] = 8'd210;
	sample_rom[112][43] = 8'd208;
	sample_rom[112][44] = 8'd203;
	sample_rom[112][45] = 8'd187;
	sample_rom[112][46] = 8'd163;
	sample_rom[112][47] = 8'd139;
	sample_rom[112][48] = 8'd116;
	sample_rom[112][49] = 8'd100;
	sample_rom[112][50] = 8'd93;
	sample_rom[112][51] = 8'd83;
	sample_rom[112][52] = 8'd68;
	sample_rom[112][53] = 8'd52;
	sample_rom[112][54] = 8'd34;
	sample_rom[112][55] = 8'd25;
	sample_rom[112][56] = 8'd27;
	sample_rom[112][57] = 8'd36;
	sample_rom[112][58] = 8'd50;
	sample_rom[112][59] = 8'd60;
	sample_rom[112][60] = 8'd65;
	sample_rom[112][61] = 8'd72;
	sample_rom[112][62] = 8'd86;
	sample_rom[112][63] = 8'd104;
	sample_rom[113][0] = 8'd130;
	sample_rom[113][1] = 8'd135;
	sample_rom[113][2] = 8'd140;
	sample_rom[113][3] = 8'd145;
	sample_rom[113][4] = 8'd149;
	sample_rom[113][5] = 8'd152;
	sample_rom[113][6] = 8'd157;
	sample_rom[113][7] = 8'd160;
	sample_rom[113][8] = 8'd164;
	sample_rom[113][9] = 8'd168;
	sample_rom[113][10] = 8'd173;
	sample_rom[113][11] = 8'd177;
	sample_rom[113][12] = 8'd180;
	sample_rom[113][13] = 8'd184;
	sample_rom[113][14] = 8'd188;
	sample_rom[113][15] = 8'd192;
	sample_rom[113][16] = 8'd195;
	sample_rom[113][17] = 8'd198;
	sample_rom[113][18] = 8'd199;
	sample_rom[113][19] = 8'd202;
	sample_rom[113][20] = 8'd204;
	sample_rom[113][21] = 8'd207;
	sample_rom[113][22] = 8'd209;
	sample_rom[113][23] = 8'd211;
	sample_rom[113][24] = 8'd213;
	sample_rom[113][25] = 8'd215;
	sample_rom[113][26] = 8'd216;
	sample_rom[113][27] = 8'd217;
	sample_rom[113][28] = 8'd218;
	sample_rom[113][29] = 8'd219;
	sample_rom[113][30] = 8'd219;
	sample_rom[113][31] = 8'd219;
	sample_rom[113][32] = 8'd219;
	sample_rom[113][33] = 8'd219;
	sample_rom[113][34] = 8'd219;
	sample_rom[113][35] = 8'd218;
	sample_rom[113][36] = 8'd217;
	sample_rom[113][37] = 8'd216;
	sample_rom[113][38] = 8'd215;
	sample_rom[113][39] = 8'd213;
	sample_rom[113][40] = 8'd211;
	sample_rom[113][41] = 8'd209;
	sample_rom[113][42] = 8'd207;
	sample_rom[113][43] = 8'd204;
	sample_rom[113][44] = 8'd202;
	sample_rom[113][45] = 8'd199;
	sample_rom[113][46] = 8'd198;
	sample_rom[113][47] = 8'd195;
	sample_rom[113][48] = 8'd192;
	sample_rom[113][49] = 8'd188;
	sample_rom[113][50] = 8'd184;
	sample_rom[113][51] = 8'd180;
	sample_rom[113][52] = 8'd177;
	sample_rom[113][53] = 8'd173;
	sample_rom[113][54] = 8'd168;
	sample_rom[113][55] = 8'd164;
	sample_rom[113][56] = 8'd160;
	sample_rom[113][57] = 8'd157;
	sample_rom[113][58] = 8'd152;
	sample_rom[113][59] = 8'd149;
	sample_rom[113][60] = 8'd145;
	sample_rom[113][61] = 8'd140;
	sample_rom[113][62] = 8'd135;
	sample_rom[113][63] = 8'd130;
	sample_rom[114][0] = 8'd131;
	sample_rom[114][1] = 8'd139;
	sample_rom[114][2] = 8'd147;
	sample_rom[114][3] = 8'd154;
	sample_rom[114][4] = 8'd160;
	sample_rom[114][5] = 8'd165;
	sample_rom[114][6] = 8'd173;
	sample_rom[114][7] = 8'd179;
	sample_rom[114][8] = 8'd185;
	sample_rom[114][9] = 8'd191;
	sample_rom[114][10] = 8'd197;
	sample_rom[114][11] = 8'd203;
	sample_rom[114][12] = 8'd207;
	sample_rom[114][13] = 8'd212;
	sample_rom[114][14] = 8'd216;
	sample_rom[114][15] = 8'd221;
	sample_rom[114][16] = 8'd223;
	sample_rom[114][17] = 8'd226;
	sample_rom[114][18] = 8'd226;
	sample_rom[114][19] = 8'd228;
	sample_rom[114][20] = 8'd229;
	sample_rom[114][21] = 8'd231;
	sample_rom[114][22] = 8'd231;
	sample_rom[114][23] = 8'd232;
	sample_rom[114][24] = 8'd232;
	sample_rom[114][25] = 8'd232;
	sample_rom[114][26] = 8'd230;
	sample_rom[114][27] = 8'd229;
	sample_rom[114][28] = 8'd227;
	sample_rom[114][29] = 8'd226;
	sample_rom[114][30] = 8'd223;
	sample_rom[114][31] = 8'd221;
	sample_rom[114][32] = 8'd218;
	sample_rom[114][33] = 8'd215;
	sample_rom[114][34] = 8'd212;
	sample_rom[114][35] = 8'd209;
	sample_rom[114][36] = 8'd206;
	sample_rom[114][37] = 8'd202;
	sample_rom[114][38] = 8'd198;
	sample_rom[114][39] = 8'd194;
	sample_rom[114][40] = 8'd190;
	sample_rom[114][41] = 8'd187;
	sample_rom[114][42] = 8'd183;
	sample_rom[114][43] = 8'd178;
	sample_rom[114][44] = 8'd175;
	sample_rom[114][45] = 8'd171;
	sample_rom[114][46] = 8'd170;
	sample_rom[114][47] = 8'd166;
	sample_rom[114][48] = 8'd163;
	sample_rom[114][49] = 8'd160;
	sample_rom[114][50] = 8'd157;
	sample_rom[114][51] = 8'd154;
	sample_rom[114][52] = 8'd152;
	sample_rom[114][53] = 8'd149;
	sample_rom[114][54] = 8'd146;
	sample_rom[114][55] = 8'd143;
	sample_rom[114][56] = 8'd141;
	sample_rom[114][57] = 8'd139;
	sample_rom[114][58] = 8'd137;
	sample_rom[114][59] = 8'd136;
	sample_rom[114][60] = 8'd135;
	sample_rom[114][61] = 8'd133;
	sample_rom[114][62] = 8'd130;
	sample_rom[114][63] = 8'd128;
	sample_rom[115][0] = 8'd131;
	sample_rom[115][1] = 8'd140;
	sample_rom[115][2] = 8'd150;
	sample_rom[115][3] = 8'd158;
	sample_rom[115][4] = 8'd166;
	sample_rom[115][5] = 8'd173;
	sample_rom[115][6] = 8'd182;
	sample_rom[115][7] = 8'd189;
	sample_rom[115][8] = 8'd195;
	sample_rom[115][9] = 8'd203;
	sample_rom[115][10] = 8'd209;
	sample_rom[115][11] = 8'd214;
	sample_rom[115][12] = 8'd220;
	sample_rom[115][13] = 8'd223;
	sample_rom[115][14] = 8'd228;
	sample_rom[115][15] = 8'd232;
	sample_rom[115][16] = 8'd234;
	sample_rom[115][17] = 8'd237;
	sample_rom[115][18] = 8'd238;
	sample_rom[115][19] = 8'd239;
	sample_rom[115][20] = 8'd238;
	sample_rom[115][21] = 8'd239;
	sample_rom[115][22] = 8'd239;
	sample_rom[115][23] = 8'd239;
	sample_rom[115][24] = 8'd236;
	sample_rom[115][25] = 8'd234;
	sample_rom[115][26] = 8'd232;
	sample_rom[115][27] = 8'd229;
	sample_rom[115][28] = 8'd225;
	sample_rom[115][29] = 8'd223;
	sample_rom[115][30] = 8'd219;
	sample_rom[115][31] = 8'd214;
	sample_rom[115][32] = 8'd210;
	sample_rom[115][33] = 8'd205;
	sample_rom[115][34] = 8'd201;
	sample_rom[115][35] = 8'd196;
	sample_rom[115][36] = 8'd191;
	sample_rom[115][37] = 8'd187;
	sample_rom[115][38] = 8'd182;
	sample_rom[115][39] = 8'd177;
	sample_rom[115][40] = 8'd173;
	sample_rom[115][41] = 8'd170;
	sample_rom[115][42] = 8'd165;
	sample_rom[115][43] = 8'd160;
	sample_rom[115][44] = 8'd157;
	sample_rom[115][45] = 8'd155;
	sample_rom[115][46] = 8'd152;
	sample_rom[115][47] = 8'd148;
	sample_rom[115][48] = 8'd145;
	sample_rom[115][49] = 8'd143;
	sample_rom[115][50] = 8'd140;
	sample_rom[115][51] = 8'd138;
	sample_rom[115][52] = 8'd136;
	sample_rom[115][53] = 8'd135;
	sample_rom[115][54] = 8'd133;
	sample_rom[115][55] = 8'd131;
	sample_rom[115][56] = 8'd130;
	sample_rom[115][57] = 8'd130;
	sample_rom[115][58] = 8'd128;
	sample_rom[115][59] = 8'd129;
	sample_rom[115][60] = 8'd128;
	sample_rom[115][61] = 8'd129;
	sample_rom[115][62] = 8'd127;
	sample_rom[115][63] = 8'd127;
	sample_rom[116][0] = 8'd131;
	sample_rom[116][1] = 8'd152;
	sample_rom[116][2] = 8'd169;
	sample_rom[116][3] = 8'd184;
	sample_rom[116][4] = 8'd199;
	sample_rom[116][5] = 8'd211;
	sample_rom[116][6] = 8'd218;
	sample_rom[116][7] = 8'd223;
	sample_rom[116][8] = 8'd224;
	sample_rom[116][9] = 8'd225;
	sample_rom[116][10] = 8'd224;
	sample_rom[116][11] = 8'd221;
	sample_rom[116][12] = 8'd219;
	sample_rom[116][13] = 8'd212;
	sample_rom[116][14] = 8'd210;
	sample_rom[116][15] = 8'd204;
	sample_rom[116][16] = 8'd199;
	sample_rom[116][17] = 8'd194;
	sample_rom[116][18] = 8'd188;
	sample_rom[116][19] = 8'd183;
	sample_rom[116][20] = 8'd179;
	sample_rom[116][21] = 8'd172;
	sample_rom[116][22] = 8'd168;
	sample_rom[116][23] = 8'd163;
	sample_rom[116][24] = 8'd161;
	sample_rom[116][25] = 8'd159;
	sample_rom[116][26] = 8'd154;
	sample_rom[116][27] = 8'd153;
	sample_rom[116][28] = 8'd152;
	sample_rom[116][29] = 8'd151;
	sample_rom[116][30] = 8'd148;
	sample_rom[116][31] = 8'd144;
	sample_rom[116][32] = 8'd143;
	sample_rom[116][33] = 8'd140;
	sample_rom[116][34] = 8'd139;
	sample_rom[116][35] = 8'd139;
	sample_rom[116][36] = 8'd138;
	sample_rom[116][37] = 8'd135;
	sample_rom[116][38] = 8'd136;
	sample_rom[116][39] = 8'd134;
	sample_rom[116][40] = 8'd136;
	sample_rom[116][41] = 8'd137;
	sample_rom[116][42] = 8'd139;
	sample_rom[116][43] = 8'd137;
	sample_rom[116][44] = 8'd139;
	sample_rom[116][45] = 8'd138;
	sample_rom[116][46] = 8'd137;
	sample_rom[116][47] = 8'd138;
	sample_rom[116][48] = 8'd137;
	sample_rom[116][49] = 8'd134;
	sample_rom[116][50] = 8'd138;
	sample_rom[116][51] = 8'd137;
	sample_rom[116][52] = 8'd135;
	sample_rom[116][53] = 8'd136;
	sample_rom[116][54] = 8'd136;
	sample_rom[116][55] = 8'd134;
	sample_rom[116][56] = 8'd136;
	sample_rom[116][57] = 8'd134;
	sample_rom[116][58] = 8'd132;
	sample_rom[116][59] = 8'd133;
	sample_rom[116][60] = 8'd132;
	sample_rom[116][61] = 8'd131;
	sample_rom[116][62] = 8'd128;
	sample_rom[116][63] = 8'd130;
	sample_rom[117][0] = 8'd131;
	sample_rom[117][1] = 8'd156;
	sample_rom[117][2] = 8'd175;
	sample_rom[117][3] = 8'd195;
	sample_rom[117][4] = 8'd211;
	sample_rom[117][5] = 8'd221;
	sample_rom[117][6] = 8'd225;
	sample_rom[117][7] = 8'd229;
	sample_rom[117][8] = 8'd225;
	sample_rom[117][9] = 8'd223;
	sample_rom[117][10] = 8'd220;
	sample_rom[117][11] = 8'd214;
	sample_rom[117][12] = 8'd209;
	sample_rom[117][13] = 8'd204;
	sample_rom[117][14] = 8'd203;
	sample_rom[117][15] = 8'd198;
	sample_rom[117][16] = 8'd195;
	sample_rom[117][17] = 8'd194;
	sample_rom[117][18] = 8'd191;
	sample_rom[117][19] = 8'd186;
	sample_rom[117][20] = 8'd185;
	sample_rom[117][21] = 8'd178;
	sample_rom[117][22] = 8'd173;
	sample_rom[117][23] = 8'd169;
	sample_rom[117][24] = 8'd164;
	sample_rom[117][25] = 8'd160;
	sample_rom[117][26] = 8'd155;
	sample_rom[117][27] = 8'd152;
	sample_rom[117][28] = 8'd148;
	sample_rom[117][29] = 8'd149;
	sample_rom[117][30] = 8'd145;
	sample_rom[117][31] = 8'd141;
	sample_rom[117][32] = 8'd141;
	sample_rom[117][33] = 8'd141;
	sample_rom[117][34] = 8'd138;
	sample_rom[117][35] = 8'd139;
	sample_rom[117][36] = 8'd139;
	sample_rom[117][37] = 8'd135;
	sample_rom[117][38] = 8'd137;
	sample_rom[117][39] = 8'd135;
	sample_rom[117][40] = 8'd136;
	sample_rom[117][41] = 8'd138;
	sample_rom[117][42] = 8'd139;
	sample_rom[117][43] = 8'd138;
	sample_rom[117][44] = 8'd139;
	sample_rom[117][45] = 8'd138;
	sample_rom[117][46] = 8'd137;
	sample_rom[117][47] = 8'd138;
	sample_rom[117][48] = 8'd137;
	sample_rom[117][49] = 8'd136;
	sample_rom[117][50] = 8'd137;
	sample_rom[117][51] = 8'd138;
	sample_rom[117][52] = 8'd136;
	sample_rom[117][53] = 8'd136;
	sample_rom[117][54] = 8'd134;
	sample_rom[117][55] = 8'd134;
	sample_rom[117][56] = 8'd136;
	sample_rom[117][57] = 8'd133;
	sample_rom[117][58] = 8'd133;
	sample_rom[117][59] = 8'd134;
	sample_rom[117][60] = 8'd131;
	sample_rom[117][61] = 8'd132;
	sample_rom[117][62] = 8'd128;
	sample_rom[117][63] = 8'd129;
	sample_rom[118][0] = 8'd132;
	sample_rom[118][1] = 8'd189;
	sample_rom[118][2] = 8'd226;
	sample_rom[118][3] = 8'd241;
	sample_rom[118][4] = 8'd234;
	sample_rom[118][5] = 8'd222;
	sample_rom[118][6] = 8'd209;
	sample_rom[118][7] = 8'd207;
	sample_rom[118][8] = 8'd203;
	sample_rom[118][9] = 8'd198;
	sample_rom[118][10] = 8'd176;
	sample_rom[118][11] = 8'd143;
	sample_rom[118][12] = 8'd107;
	sample_rom[118][13] = 8'd71;
	sample_rom[118][14] = 8'd53;
	sample_rom[118][15] = 8'd51;
	sample_rom[118][16] = 8'd64;
	sample_rom[118][17] = 8'd88;
	sample_rom[118][18] = 8'd104;
	sample_rom[118][19] = 8'd112;
	sample_rom[118][20] = 8'd112;
	sample_rom[118][21] = 8'd105;
	sample_rom[118][22] = 8'd106;
	sample_rom[118][23] = 8'd110;
	sample_rom[118][24] = 8'd123;
	sample_rom[118][25] = 8'd138;
	sample_rom[118][26] = 8'd145;
	sample_rom[118][27] = 8'd147;
	sample_rom[118][28] = 8'd135;
	sample_rom[118][29] = 8'd124;
	sample_rom[118][30] = 8'd113;
	sample_rom[118][31] = 8'd116;
	sample_rom[118][32] = 8'd123;
	sample_rom[118][33] = 8'd135;
	sample_rom[118][34] = 8'd148;
	sample_rom[118][35] = 8'd157;
	sample_rom[118][36] = 8'd157;
	sample_rom[118][37] = 8'd153;
	sample_rom[118][38] = 8'd147;
	sample_rom[118][39] = 8'd142;
	sample_rom[118][40] = 8'd142;
	sample_rom[118][41] = 8'd143;
	sample_rom[118][42] = 8'd142;
	sample_rom[118][43] = 8'd143;
	sample_rom[118][44] = 8'd136;
	sample_rom[118][45] = 8'd125;
	sample_rom[118][46] = 8'd114;
	sample_rom[118][47] = 8'd104;
	sample_rom[118][48] = 8'd101;
	sample_rom[118][49] = 8'd104;
	sample_rom[118][50] = 8'd109;
	sample_rom[118][51] = 8'd114;
	sample_rom[118][52] = 8'd121;
	sample_rom[118][53] = 8'd122;
	sample_rom[118][54] = 8'd123;
	sample_rom[118][55] = 8'd122;
	sample_rom[118][56] = 8'd126;
	sample_rom[118][57] = 8'd127;
	sample_rom[118][58] = 8'd127;
	sample_rom[118][59] = 8'd130;
	sample_rom[118][60] = 8'd132;
	sample_rom[118][61] = 8'd135;
	sample_rom[118][62] = 8'd137;
	sample_rom[118][63] = 8'd133;
	sample_rom[119][0] = 8'd132;
	sample_rom[119][1] = 8'd197;
	sample_rom[119][2] = 8'd240;
	sample_rom[119][3] = 8'd249;
	sample_rom[119][4] = 8'd234;
	sample_rom[119][5] = 8'd212;
	sample_rom[119][6] = 8'd202;
	sample_rom[119][7] = 8'd206;
	sample_rom[119][8] = 8'd222;
	sample_rom[119][9] = 8'd230;
	sample_rom[119][10] = 8'd221;
	sample_rom[119][11] = 8'd188;
	sample_rom[119][12] = 8'd142;
	sample_rom[119][13] = 8'd96;
	sample_rom[119][14] = 8'd65;
	sample_rom[119][15] = 8'd54;
	sample_rom[119][16] = 8'd62;
	sample_rom[119][17] = 8'd82;
	sample_rom[119][18] = 8'd101;
	sample_rom[119][19] = 8'd109;
	sample_rom[119][20] = 8'd108;
	sample_rom[119][21] = 8'd97;
	sample_rom[119][22] = 8'd92;
	sample_rom[119][23] = 8'd93;
	sample_rom[119][24] = 8'd106;
	sample_rom[119][25] = 8'd128;
	sample_rom[119][26] = 8'd149;
	sample_rom[119][27] = 8'd154;
	sample_rom[119][28] = 8'd143;
	sample_rom[119][29] = 8'd127;
	sample_rom[119][30] = 8'd113;
	sample_rom[119][31] = 8'd103;
	sample_rom[119][32] = 8'd107;
	sample_rom[119][33] = 8'd119;
	sample_rom[119][34] = 8'd132;
	sample_rom[119][35] = 8'd144;
	sample_rom[119][36] = 8'd150;
	sample_rom[119][37] = 8'd151;
	sample_rom[119][38] = 8'd148;
	sample_rom[119][39] = 8'd148;
	sample_rom[119][40] = 8'd150;
	sample_rom[119][41] = 8'd156;
	sample_rom[119][42] = 8'd163;
	sample_rom[119][43] = 8'd167;
	sample_rom[119][44] = 8'd165;
	sample_rom[119][45] = 8'd157;
	sample_rom[119][46] = 8'd143;
	sample_rom[119][47] = 8'd129;
	sample_rom[119][48] = 8'd116;
	sample_rom[119][49] = 8'd113;
	sample_rom[119][50] = 8'd110;
	sample_rom[119][51] = 8'd111;
	sample_rom[119][52] = 8'd111;
	sample_rom[119][53] = 8'd113;
	sample_rom[119][54] = 8'd112;
	sample_rom[119][55] = 8'd113;
	sample_rom[119][56] = 8'd114;
	sample_rom[119][57] = 8'd118;
	sample_rom[119][58] = 8'd122;
	sample_rom[119][59] = 8'd129;
	sample_rom[119][60] = 8'd131;
	sample_rom[119][61] = 8'd138;
	sample_rom[119][62] = 8'd138;
	sample_rom[119][63] = 8'd133;
	sample_rom[120][0] = 8'd128;
	sample_rom[120][1] = 8'd196;
	sample_rom[120][2] = 8'd229;
	sample_rom[120][3] = 8'd225;
	sample_rom[120][4] = 8'd198;
	sample_rom[120][5] = 8'd168;
	sample_rom[120][6] = 8'd152;
	sample_rom[120][7] = 8'd159;
	sample_rom[120][8] = 8'd173;
	sample_rom[120][9] = 8'd195;
	sample_rom[120][10] = 8'd208;
	sample_rom[120][11] = 8'd200;
	sample_rom[120][12] = 8'd174;
	sample_rom[120][13] = 8'd136;
	sample_rom[120][14] = 8'd103;
	sample_rom[120][15] = 8'd85;
	sample_rom[120][16] = 8'd77;
	sample_rom[120][17] = 8'd88;
	sample_rom[120][18] = 8'd101;
	sample_rom[120][19] = 8'd113;
	sample_rom[120][20] = 8'd120;
	sample_rom[120][21] = 8'd118;
	sample_rom[120][22] = 8'd114;
	sample_rom[120][23] = 8'd111;
	sample_rom[120][24] = 8'd112;
	sample_rom[120][25] = 8'd123;
	sample_rom[120][26] = 8'd126;
	sample_rom[120][27] = 8'd135;
	sample_rom[120][28] = 8'd139;
	sample_rom[120][29] = 8'd144;
	sample_rom[120][30] = 8'd143;
	sample_rom[120][31] = 8'd140;
	sample_rom[120][32] = 8'd135;
	sample_rom[120][33] = 8'd133;
	sample_rom[120][34] = 8'd131;
	sample_rom[120][35] = 8'd127;
	sample_rom[120][36] = 8'd124;
	sample_rom[120][37] = 8'd121;
	sample_rom[120][38] = 8'd123;
	sample_rom[120][39] = 8'd128;
	sample_rom[120][40] = 8'd135;
	sample_rom[120][41] = 8'd143;
	sample_rom[120][42] = 8'd147;
	sample_rom[120][43] = 8'd149;
	sample_rom[120][44] = 8'd146;
	sample_rom[120][45] = 8'd143;
	sample_rom[120][46] = 8'd141;
	sample_rom[120][47] = 8'd142;
	sample_rom[120][48] = 8'd143;
	sample_rom[120][49] = 8'd143;
	sample_rom[120][50] = 8'd142;
	sample_rom[120][51] = 8'd146;
	sample_rom[120][52] = 8'd148;
	sample_rom[120][53] = 8'd139;
	sample_rom[120][54] = 8'd132;
	sample_rom[120][55] = 8'd123;
	sample_rom[120][56] = 8'd121;
	sample_rom[120][57] = 8'd122;
	sample_rom[120][58] = 8'd122;
	sample_rom[120][59] = 8'd125;
	sample_rom[120][60] = 8'd126;
	sample_rom[120][61] = 8'd131;
	sample_rom[120][62] = 8'd135;
	sample_rom[120][63] = 8'd133;
	sample_rom[121][0] = 8'd128;
	sample_rom[121][1] = 8'd195;
	sample_rom[121][2] = 8'd231;
	sample_rom[121][3] = 8'd230;
	sample_rom[121][4] = 8'd202;
	sample_rom[121][5] = 8'd162;
	sample_rom[121][6] = 8'd124;
	sample_rom[121][7] = 8'd110;
	sample_rom[121][8] = 8'd112;
	sample_rom[121][9] = 8'd134;
	sample_rom[121][10] = 8'd161;
	sample_rom[121][11] = 8'd184;
	sample_rom[121][12] = 8'd197;
	sample_rom[121][13] = 8'd193;
	sample_rom[121][14] = 8'd173;
	sample_rom[121][15] = 8'd143;
	sample_rom[121][16] = 8'd117;
	sample_rom[121][17] = 8'd100;
	sample_rom[121][18] = 8'd95;
	sample_rom[121][19] = 8'd96;
	sample_rom[121][20] = 8'd100;
	sample_rom[121][21] = 8'd109;
	sample_rom[121][22] = 8'd114;
	sample_rom[121][23] = 8'd114;
	sample_rom[121][24] = 8'd113;
	sample_rom[121][25] = 8'd114;
	sample_rom[121][26] = 8'd117;
	sample_rom[121][27] = 8'd118;
	sample_rom[121][28] = 8'd125;
	sample_rom[121][29] = 8'd128;
	sample_rom[121][30] = 8'd131;
	sample_rom[121][31] = 8'd132;
	sample_rom[121][32] = 8'd130;
	sample_rom[121][33] = 8'd128;
	sample_rom[121][34] = 8'd133;
	sample_rom[121][35] = 8'd137;
	sample_rom[121][36] = 8'd144;
	sample_rom[121][37] = 8'd145;
	sample_rom[121][38] = 8'd148;
	sample_rom[121][39] = 8'd143;
	sample_rom[121][40] = 8'd136;
	sample_rom[121][41] = 8'd126;
	sample_rom[121][42] = 8'd124;
	sample_rom[121][43] = 8'd127;
	sample_rom[121][44] = 8'd128;
	sample_rom[121][45] = 8'd129;
	sample_rom[121][46] = 8'd128;
	sample_rom[121][47] = 8'd128;
	sample_rom[121][48] = 8'd130;
	sample_rom[121][49] = 8'd129;
	sample_rom[121][50] = 8'd134;
	sample_rom[121][51] = 8'd138;
	sample_rom[121][52] = 8'd141;
	sample_rom[121][53] = 8'd145;
	sample_rom[121][54] = 8'd146;
	sample_rom[121][55] = 8'd146;
	sample_rom[121][56] = 8'd146;
	sample_rom[121][57] = 8'd142;
	sample_rom[121][58] = 8'd139;
	sample_rom[121][59] = 8'd141;
	sample_rom[121][60] = 8'd145;
	sample_rom[121][61] = 8'd141;
	sample_rom[121][62] = 8'd135;
	sample_rom[121][63] = 8'd131;
	sample_rom[122][0] = 8'd128;
	sample_rom[122][1] = 8'd194;
	sample_rom[122][2] = 8'd233;
	sample_rom[122][3] = 8'd237;
	sample_rom[122][4] = 8'd216;
	sample_rom[122][5] = 8'd181;
	sample_rom[122][6] = 8'd140;
	sample_rom[122][7] = 8'd113;
	sample_rom[122][8] = 8'd104;
	sample_rom[122][9] = 8'd111;
	sample_rom[122][10] = 8'd136;
	sample_rom[122][11] = 8'd162;
	sample_rom[122][12] = 8'd190;
	sample_rom[122][13] = 8'd202;
	sample_rom[122][14] = 8'd201;
	sample_rom[122][15] = 8'd188;
	sample_rom[122][16] = 8'd167;
	sample_rom[122][17] = 8'd144;
	sample_rom[122][18] = 8'd127;
	sample_rom[122][19] = 8'd119;
	sample_rom[122][20] = 8'd120;
	sample_rom[122][21] = 8'd125;
	sample_rom[122][22] = 8'd134;
	sample_rom[122][23] = 8'd139;
	sample_rom[122][24] = 8'd145;
	sample_rom[122][25] = 8'd143;
	sample_rom[122][26] = 8'd137;
	sample_rom[122][27] = 8'd126;
	sample_rom[122][28] = 8'd119;
	sample_rom[122][29] = 8'd110;
	sample_rom[122][30] = 8'd109;
	sample_rom[122][31] = 8'd109;
	sample_rom[122][32] = 8'd115;
	sample_rom[122][33] = 8'd116;
	sample_rom[122][34] = 8'd116;
	sample_rom[122][35] = 8'd116;
	sample_rom[122][36] = 8'd113;
	sample_rom[122][37] = 8'd114;
	sample_rom[122][38] = 8'd111;
	sample_rom[122][39] = 8'd112;
	sample_rom[122][40] = 8'd116;
	sample_rom[122][41] = 8'd123;
	sample_rom[122][42] = 8'd126;
	sample_rom[122][43] = 8'd127;
	sample_rom[122][44] = 8'd130;
	sample_rom[122][45] = 8'd129;
	sample_rom[122][46] = 8'd123;
	sample_rom[122][47] = 8'd122;
	sample_rom[122][48] = 8'd121;
	sample_rom[122][49] = 8'd118;
	sample_rom[122][50] = 8'd122;
	sample_rom[122][51] = 8'd132;
	sample_rom[122][52] = 8'd137;
	sample_rom[122][53] = 8'd135;
	sample_rom[122][54] = 8'd133;
	sample_rom[122][55] = 8'd131;
	sample_rom[122][56] = 8'd129;
	sample_rom[122][57] = 8'd126;
	sample_rom[122][58] = 8'd126;
	sample_rom[122][59] = 8'd125;
	sample_rom[122][60] = 8'd129;
	sample_rom[122][61] = 8'd132;
	sample_rom[122][62] = 8'd136;
	sample_rom[122][63] = 8'd133;
	sample_rom[123][0] = 8'd133;
	sample_rom[123][1] = 8'd183;
	sample_rom[123][2] = 8'd219;
	sample_rom[123][3] = 8'd239;
	sample_rom[123][4] = 8'd238;
	sample_rom[123][5] = 8'd219;
	sample_rom[123][6] = 8'd188;
	sample_rom[123][7] = 8'd154;
	sample_rom[123][8] = 8'd125;
	sample_rom[123][9] = 8'd106;
	sample_rom[123][10] = 8'd105;
	sample_rom[123][11] = 8'd116;
	sample_rom[123][12] = 8'd138;
	sample_rom[123][13] = 8'd164;
	sample_rom[123][14] = 8'd189;
	sample_rom[123][15] = 8'd211;
	sample_rom[123][16] = 8'd220;
	sample_rom[123][17] = 8'd220;
	sample_rom[123][18] = 8'd207;
	sample_rom[123][19] = 8'd188;
	sample_rom[123][20] = 8'd161;
	sample_rom[123][21] = 8'd138;
	sample_rom[123][22] = 8'd119;
	sample_rom[123][23] = 8'd107;
	sample_rom[123][24] = 8'd106;
	sample_rom[123][25] = 8'd107;
	sample_rom[123][26] = 8'd110;
	sample_rom[123][27] = 8'd116;
	sample_rom[123][28] = 8'd118;
	sample_rom[123][29] = 8'd117;
	sample_rom[123][30] = 8'd113;
	sample_rom[123][31] = 8'd110;
	sample_rom[123][32] = 8'd104;
	sample_rom[123][33] = 8'd100;
	sample_rom[123][34] = 8'd99;
	sample_rom[123][35] = 8'd99;
	sample_rom[123][36] = 8'd100;
	sample_rom[123][37] = 8'd98;
	sample_rom[123][38] = 8'd100;
	sample_rom[123][39] = 8'd100;
	sample_rom[123][40] = 8'd102;
	sample_rom[123][41] = 8'd101;
	sample_rom[123][42] = 8'd100;
	sample_rom[123][43] = 8'd103;
	sample_rom[123][44] = 8'd103;
	sample_rom[123][45] = 8'd106;
	sample_rom[123][46] = 8'd113;
	sample_rom[123][47] = 8'd119;
	sample_rom[123][48] = 8'd127;
	sample_rom[123][49] = 8'd134;
	sample_rom[123][50] = 8'd141;
	sample_rom[123][51] = 8'd142;
	sample_rom[123][52] = 8'd143;
	sample_rom[123][53] = 8'd143;
	sample_rom[123][54] = 8'd140;
	sample_rom[123][55] = 8'd137;
	sample_rom[123][56] = 8'd136;
	sample_rom[123][57] = 8'd134;
	sample_rom[123][58] = 8'd131;
	sample_rom[123][59] = 8'd128;
	sample_rom[123][60] = 8'd128;
	sample_rom[123][61] = 8'd128;
	sample_rom[123][62] = 8'd129;
	sample_rom[123][63] = 8'd129;
	sample_rom[124][0] = 8'd131;
	sample_rom[124][1] = 8'd160;
	sample_rom[124][2] = 8'd186;
	sample_rom[124][3] = 8'd207;
	sample_rom[124][4] = 8'd218;
	sample_rom[124][5] = 8'd223;
	sample_rom[124][6] = 8'd221;
	sample_rom[124][7] = 8'd207;
	sample_rom[124][8] = 8'd187;
	sample_rom[124][9] = 8'd165;
	sample_rom[124][10] = 8'd142;
	sample_rom[124][11] = 8'd121;
	sample_rom[124][12] = 8'd105;
	sample_rom[124][13] = 8'd95;
	sample_rom[124][14] = 8'd92;
	sample_rom[124][15] = 8'd97;
	sample_rom[124][16] = 8'd104;
	sample_rom[124][17] = 8'd121;
	sample_rom[124][18] = 8'd138;
	sample_rom[124][19] = 8'd156;
	sample_rom[124][20] = 8'd174;
	sample_rom[124][21] = 8'd189;
	sample_rom[124][22] = 8'd200;
	sample_rom[124][23] = 8'd202;
	sample_rom[124][24] = 8'd200;
	sample_rom[124][25] = 8'd191;
	sample_rom[124][26] = 8'd179;
	sample_rom[124][27] = 8'd165;
	sample_rom[124][28] = 8'd147;
	sample_rom[124][29] = 8'd129;
	sample_rom[124][30] = 8'd114;
	sample_rom[124][31] = 8'd101;
	sample_rom[124][32] = 8'd93;
	sample_rom[124][33] = 8'd87;
	sample_rom[124][34] = 8'd85;
	sample_rom[124][35] = 8'd86;
	sample_rom[124][36] = 8'd91;
	sample_rom[124][37] = 8'd96;
	sample_rom[124][38] = 8'd102;
	sample_rom[124][39] = 8'd106;
	sample_rom[124][40] = 8'd113;
	sample_rom[124][41] = 8'd118;
	sample_rom[124][42] = 8'd121;
	sample_rom[124][43] = 8'd122;
	sample_rom[124][44] = 8'd121;
	sample_rom[124][45] = 8'd118;
	sample_rom[124][46] = 8'd115;
	sample_rom[124][47] = 8'd112;
	sample_rom[124][48] = 8'd107;
	sample_rom[124][49] = 8'd103;
	sample_rom[124][50] = 8'd101;
	sample_rom[124][51] = 8'd98;
	sample_rom[124][52] = 8'd97;
	sample_rom[124][53] = 8'd97;
	sample_rom[124][54] = 8'd97;
	sample_rom[124][55] = 8'd98;
	sample_rom[124][56] = 8'd101;
	sample_rom[124][57] = 8'd106;
	sample_rom[124][58] = 8'd109;
	sample_rom[124][59] = 8'd112;
	sample_rom[124][60] = 8'd116;
	sample_rom[124][61] = 8'd119;
	sample_rom[124][62] = 8'd123;
	sample_rom[124][63] = 8'd126;
	sample_rom[125][0] = 8'd132;
	sample_rom[125][1] = 8'd156;
	sample_rom[125][2] = 8'd179;
	sample_rom[125][3] = 8'd199;
	sample_rom[125][4] = 8'd214;
	sample_rom[125][5] = 8'd225;
	sample_rom[125][6] = 8'd229;
	sample_rom[125][7] = 8'd227;
	sample_rom[125][8] = 8'd222;
	sample_rom[125][9] = 8'd209;
	sample_rom[125][10] = 8'd196;
	sample_rom[125][11] = 8'd177;
	sample_rom[125][12] = 8'd160;
	sample_rom[125][13] = 8'd144;
	sample_rom[125][14] = 8'd129;
	sample_rom[125][15] = 8'd117;
	sample_rom[125][16] = 8'd110;
	sample_rom[125][17] = 8'd108;
	sample_rom[125][18] = 8'd109;
	sample_rom[125][19] = 8'd116;
	sample_rom[125][20] = 8'd127;
	sample_rom[125][21] = 8'd139;
	sample_rom[125][22] = 8'd155;
	sample_rom[125][23] = 8'd170;
	sample_rom[125][24] = 8'd186;
	sample_rom[125][25] = 8'd197;
	sample_rom[125][26] = 8'd209;
	sample_rom[125][27] = 8'd215;
	sample_rom[125][28] = 8'd219;
	sample_rom[125][29] = 8'd218;
	sample_rom[125][30] = 8'd213;
	sample_rom[125][31] = 8'd204;
	sample_rom[125][32] = 8'd190;
	sample_rom[125][33] = 8'd177;
	sample_rom[125][34] = 8'd162;
	sample_rom[125][35] = 8'd148;
	sample_rom[125][36] = 8'd133;
	sample_rom[125][37] = 8'd120;
	sample_rom[125][38] = 8'd109;
	sample_rom[125][39] = 8'd101;
	sample_rom[125][40] = 8'd97;
	sample_rom[125][41] = 8'd97;
	sample_rom[125][42] = 8'd97;
	sample_rom[125][43] = 8'd102;
	sample_rom[125][44] = 8'd105;
	sample_rom[125][45] = 8'd112;
	sample_rom[125][46] = 8'd119;
	sample_rom[125][47] = 8'd124;
	sample_rom[125][48] = 8'd130;
	sample_rom[125][49] = 8'd134;
	sample_rom[125][50] = 8'd137;
	sample_rom[125][51] = 8'd138;
	sample_rom[125][52] = 8'd138;
	sample_rom[125][53] = 8'd136;
	sample_rom[125][54] = 8'd134;
	sample_rom[125][55] = 8'd130;
	sample_rom[125][56] = 8'd127;
	sample_rom[125][57] = 8'd125;
	sample_rom[125][58] = 8'd124;
	sample_rom[125][59] = 8'd123;
	sample_rom[125][60] = 8'd122;
	sample_rom[125][61] = 8'd123;
	sample_rom[125][62] = 8'd122;
	sample_rom[125][63] = 8'd128;
	sample_rom[126][0] = 8'd131;
	sample_rom[126][1] = 8'd148;
	sample_rom[126][2] = 8'd161;
	sample_rom[126][3] = 8'd177;
	sample_rom[126][4] = 8'd187;
	sample_rom[126][5] = 8'd196;
	sample_rom[126][6] = 8'd202;
	sample_rom[126][7] = 8'd204;
	sample_rom[126][8] = 8'd204;
	sample_rom[126][9] = 8'd199;
	sample_rom[126][10] = 8'd192;
	sample_rom[126][11] = 8'd184;
	sample_rom[126][12] = 8'd173;
	sample_rom[126][13] = 8'd161;
	sample_rom[126][14] = 8'd149;
	sample_rom[126][15] = 8'd138;
	sample_rom[126][16] = 8'd127;
	sample_rom[126][17] = 8'd117;
	sample_rom[126][18] = 8'd111;
	sample_rom[126][19] = 8'd105;
	sample_rom[126][20] = 8'd103;
	sample_rom[126][21] = 8'd105;
	sample_rom[126][22] = 8'd107;
	sample_rom[126][23] = 8'd114;
	sample_rom[126][24] = 8'd122;
	sample_rom[126][25] = 8'd133;
	sample_rom[126][26] = 8'd144;
	sample_rom[126][27] = 8'd155;
	sample_rom[126][28] = 8'd165;
	sample_rom[126][29] = 8'd175;
	sample_rom[126][30] = 8'd186;
	sample_rom[126][31] = 8'd194;
	sample_rom[126][32] = 8'd200;
	sample_rom[126][33] = 8'd203;
	sample_rom[126][34] = 8'd203;
	sample_rom[126][35] = 8'd204;
	sample_rom[126][36] = 8'd201;
	sample_rom[126][37] = 8'd195;
	sample_rom[126][38] = 8'd190;
	sample_rom[126][39] = 8'd181;
	sample_rom[126][40] = 8'd174;
	sample_rom[126][41] = 8'd165;
	sample_rom[126][42] = 8'd159;
	sample_rom[126][43] = 8'd151;
	sample_rom[126][44] = 8'd145;
	sample_rom[126][45] = 8'd138;
	sample_rom[126][46] = 8'd135;
	sample_rom[126][47] = 8'd133;
	sample_rom[126][48] = 8'd131;
	sample_rom[126][49] = 8'd130;
	sample_rom[126][50] = 8'd133;
	sample_rom[126][51] = 8'd132;
	sample_rom[126][52] = 8'd136;
	sample_rom[126][53] = 8'd137;
	sample_rom[126][54] = 8'd140;
	sample_rom[126][55] = 8'd142;
	sample_rom[126][56] = 8'd143;
	sample_rom[126][57] = 8'd143;
	sample_rom[126][58] = 8'd144;
	sample_rom[126][59] = 8'd143;
	sample_rom[126][60] = 8'd141;
	sample_rom[126][61] = 8'd140;
	sample_rom[126][62] = 8'd135;
	sample_rom[126][63] = 8'd132;
	sample_rom[127][0] = 8'd131;
	sample_rom[127][1] = 8'd141;
	sample_rom[127][2] = 8'd151;
	sample_rom[127][3] = 8'd160;
	sample_rom[127][4] = 8'd168;
	sample_rom[127][5] = 8'd175;
	sample_rom[127][6] = 8'd181;
	sample_rom[127][7] = 8'd187;
	sample_rom[127][8] = 8'd190;
	sample_rom[127][9] = 8'd193;
	sample_rom[127][10] = 8'd194;
	sample_rom[127][11] = 8'd193;
	sample_rom[127][12] = 8'd191;
	sample_rom[127][13] = 8'd187;
	sample_rom[127][14] = 8'd184;
	sample_rom[127][15] = 8'd179;
	sample_rom[127][16] = 8'd173;
	sample_rom[127][17] = 8'd166;
	sample_rom[127][18] = 8'd160;
	sample_rom[127][19] = 8'd155;
	sample_rom[127][20] = 8'd149;
	sample_rom[127][21] = 8'd145;
	sample_rom[127][22] = 8'd139;
	sample_rom[127][23] = 8'd136;
	sample_rom[127][24] = 8'd133;
	sample_rom[127][25] = 8'd132;
	sample_rom[127][26] = 8'd131;
	sample_rom[127][27] = 8'd132;
	sample_rom[127][28] = 8'd134;
	sample_rom[127][29] = 8'd136;
	sample_rom[127][30] = 8'd139;
	sample_rom[127][31] = 8'd143;
	sample_rom[127][32] = 8'd148;
	sample_rom[127][33] = 8'd153;
	sample_rom[127][34] = 8'd158;
	sample_rom[127][35] = 8'd163;
	sample_rom[127][36] = 8'd167;
	sample_rom[127][37] = 8'd172;
	sample_rom[127][38] = 8'd176;
	sample_rom[127][39] = 8'd180;
	sample_rom[127][40] = 8'd183;
	sample_rom[127][41] = 8'd183;
	sample_rom[127][42] = 8'd185;
	sample_rom[127][43] = 8'd184;
	sample_rom[127][44] = 8'd183;
	sample_rom[127][45] = 8'd181;
	sample_rom[127][46] = 8'd179;
	sample_rom[127][47] = 8'd176;
	sample_rom[127][48] = 8'd173;
	sample_rom[127][49] = 8'd168;
	sample_rom[127][50] = 8'd163;
	sample_rom[127][51] = 8'd160;
	sample_rom[127][52] = 8'd156;
	sample_rom[127][53] = 8'd151;
	sample_rom[127][54] = 8'd147;
	sample_rom[127][55] = 8'd142;
	sample_rom[127][56] = 8'd139;
	sample_rom[127][57] = 8'd136;
	sample_rom[127][58] = 8'd134;
	sample_rom[127][59] = 8'd133;
	sample_rom[127][60] = 8'd131;
	sample_rom[127][61] = 8'd130;
	sample_rom[127][62] = 8'd128;
	sample_rom[127][63] = 8'd128;
	sample_rom[128][0] = 8'd130;
	sample_rom[128][1] = 8'd138;
	sample_rom[128][2] = 8'd146;
	sample_rom[128][3] = 8'd154;
	sample_rom[128][4] = 8'd160;
	sample_rom[128][5] = 8'd168;
	sample_rom[128][6] = 8'd173;
	sample_rom[128][7] = 8'd179;
	sample_rom[128][8] = 8'd183;
	sample_rom[128][9] = 8'd187;
	sample_rom[128][10] = 8'd189;
	sample_rom[128][11] = 8'd192;
	sample_rom[128][12] = 8'd192;
	sample_rom[128][13] = 8'd191;
	sample_rom[128][14] = 8'd192;
	sample_rom[128][15] = 8'd190;
	sample_rom[128][16] = 8'd187;
	sample_rom[128][17] = 8'd183;
	sample_rom[128][18] = 8'd179;
	sample_rom[128][19] = 8'd173;
	sample_rom[128][20] = 8'd168;
	sample_rom[128][21] = 8'd163;
	sample_rom[128][22] = 8'd158;
	sample_rom[128][23] = 8'd154;
	sample_rom[128][24] = 8'd147;
	sample_rom[128][25] = 8'd142;
	sample_rom[128][26] = 8'd136;
	sample_rom[128][27] = 8'd132;
	sample_rom[128][28] = 8'd129;
	sample_rom[128][29] = 8'd125;
	sample_rom[128][30] = 8'd123;
	sample_rom[128][31] = 8'd122;
	sample_rom[128][32] = 8'd121;
	sample_rom[128][33] = 8'd120;
	sample_rom[128][34] = 8'd120;
	sample_rom[128][35] = 8'd122;
	sample_rom[128][36] = 8'd124;
	sample_rom[128][37] = 8'd125;
	sample_rom[128][38] = 8'd130;
	sample_rom[128][39] = 8'd133;
	sample_rom[128][40] = 8'd138;
	sample_rom[128][41] = 8'd142;
	sample_rom[128][42] = 8'd147;
	sample_rom[128][43] = 8'd151;
	sample_rom[128][44] = 8'd157;
	sample_rom[128][45] = 8'd160;
	sample_rom[128][46] = 8'd164;
	sample_rom[128][47] = 8'd168;
	sample_rom[128][48] = 8'd172;
	sample_rom[128][49] = 8'd174;
	sample_rom[128][50] = 8'd176;
	sample_rom[128][51] = 8'd177;
	sample_rom[128][52] = 8'd178;
	sample_rom[128][53] = 8'd176;
	sample_rom[128][54] = 8'd176;
	sample_rom[128][55] = 8'd173;
	sample_rom[128][56] = 8'd171;
	sample_rom[128][57] = 8'd166;
	sample_rom[128][58] = 8'd163;
	sample_rom[128][59] = 8'd159;
	sample_rom[128][60] = 8'd153;
	sample_rom[128][61] = 8'd146;
	sample_rom[128][62] = 8'd140;
	sample_rom[128][63] = 8'd133;
	sample_rom[129][0] = 8'd129;
	sample_rom[129][1] = 8'd133;
	sample_rom[129][2] = 8'd137;
	sample_rom[129][3] = 8'd140;
	sample_rom[129][4] = 8'd143;
	sample_rom[129][5] = 8'd147;
	sample_rom[129][6] = 8'd150;
	sample_rom[129][7] = 8'd153;
	sample_rom[129][8] = 8'd156;
	sample_rom[129][9] = 8'd158;
	sample_rom[129][10] = 8'd160;
	sample_rom[129][11] = 8'd161;
	sample_rom[129][12] = 8'd163;
	sample_rom[129][13] = 8'd164;
	sample_rom[129][14] = 8'd165;
	sample_rom[129][15] = 8'd165;
	sample_rom[129][16] = 8'd165;
	sample_rom[129][17] = 8'd165;
	sample_rom[129][18] = 8'd165;
	sample_rom[129][19] = 8'd164;
	sample_rom[129][20] = 8'd162;
	sample_rom[129][21] = 8'd160;
	sample_rom[129][22] = 8'd159;
	sample_rom[129][23] = 8'd157;
	sample_rom[129][24] = 8'd155;
	sample_rom[129][25] = 8'd152;
	sample_rom[129][26] = 8'd149;
	sample_rom[129][27] = 8'd145;
	sample_rom[129][28] = 8'd142;
	sample_rom[129][29] = 8'd138;
	sample_rom[129][30] = 8'd135;
	sample_rom[129][31] = 8'd131;
	sample_rom[129][32] = 8'd127;
	sample_rom[129][33] = 8'd123;
	sample_rom[129][34] = 8'd119;
	sample_rom[129][35] = 8'd116;
	sample_rom[129][36] = 8'd113;
	sample_rom[129][37] = 8'd109;
	sample_rom[129][38] = 8'd106;
	sample_rom[129][39] = 8'd103;
	sample_rom[129][40] = 8'd100;
	sample_rom[129][41] = 8'd98;
	sample_rom[129][42] = 8'd97;
	sample_rom[129][43] = 8'd95;
	sample_rom[129][44] = 8'd93;
	sample_rom[129][45] = 8'd92;
	sample_rom[129][46] = 8'd91;
	sample_rom[129][47] = 8'd91;
	sample_rom[129][48] = 8'd91;
	sample_rom[129][49] = 8'd91;
	sample_rom[129][50] = 8'd92;
	sample_rom[129][51] = 8'd92;
	sample_rom[129][52] = 8'd94;
	sample_rom[129][53] = 8'd96;
	sample_rom[129][54] = 8'd97;
	sample_rom[129][55] = 8'd99;
	sample_rom[129][56] = 8'd101;
	sample_rom[129][57] = 8'd104;
	sample_rom[129][58] = 8'd107;
	sample_rom[129][59] = 8'd111;
	sample_rom[129][60] = 8'd114;
	sample_rom[129][61] = 8'd118;
	sample_rom[129][62] = 8'd121;
	sample_rom[129][63] = 8'd125;
	sample_rom[130][0] = 8'd130;
	sample_rom[130][1] = 8'd200;
	sample_rom[130][2] = 8'd227;
	sample_rom[130][3] = 8'd223;
	sample_rom[130][4] = 8'd211;
	sample_rom[130][5] = 8'd214;
	sample_rom[130][6] = 8'd219;
	sample_rom[130][7] = 8'd222;
	sample_rom[130][8] = 8'd220;
	sample_rom[130][9] = 8'd223;
	sample_rom[130][10] = 8'd231;
	sample_rom[130][11] = 8'd236;
	sample_rom[130][12] = 8'd231;
	sample_rom[130][13] = 8'd219;
	sample_rom[130][14] = 8'd210;
	sample_rom[130][15] = 8'd204;
	sample_rom[130][16] = 8'd197;
	sample_rom[130][17] = 8'd190;
	sample_rom[130][18] = 8'd184;
	sample_rom[130][19] = 8'd183;
	sample_rom[130][20] = 8'd184;
	sample_rom[130][21] = 8'd175;
	sample_rom[130][22] = 8'd166;
	sample_rom[130][23] = 8'd160;
	sample_rom[130][24] = 8'd159;
	sample_rom[130][25] = 8'd153;
	sample_rom[130][26] = 8'd149;
	sample_rom[130][27] = 8'd148;
	sample_rom[130][28] = 8'd142;
	sample_rom[130][29] = 8'd144;
	sample_rom[130][30] = 8'd139;
	sample_rom[130][31] = 8'd131;
	sample_rom[130][32] = 8'd125;
	sample_rom[130][33] = 8'd126;
	sample_rom[130][34] = 8'd121;
	sample_rom[130][35] = 8'd117;
	sample_rom[130][36] = 8'd118;
	sample_rom[130][37] = 8'd116;
	sample_rom[130][38] = 8'd118;
	sample_rom[130][39] = 8'd115;
	sample_rom[130][40] = 8'd113;
	sample_rom[130][41] = 8'd114;
	sample_rom[130][42] = 8'd120;
	sample_rom[130][43] = 8'd121;
	sample_rom[130][44] = 8'd125;
	sample_rom[130][45] = 8'd125;
	sample_rom[130][46] = 8'd128;
	sample_rom[130][47] = 8'd134;
	sample_rom[130][48] = 8'd133;
	sample_rom[130][49] = 8'd132;
	sample_rom[130][50] = 8'd132;
	sample_rom[130][51] = 8'd133;
	sample_rom[130][52] = 8'd139;
	sample_rom[130][53] = 8'd137;
	sample_rom[130][54] = 8'd139;
	sample_rom[130][55] = 8'd138;
	sample_rom[130][56] = 8'd138;
	sample_rom[130][57] = 8'd133;
	sample_rom[130][58] = 8'd136;
	sample_rom[130][59] = 8'd136;
	sample_rom[130][60] = 8'd132;
	sample_rom[130][61] = 8'd137;
	sample_rom[130][62] = 8'd129;
	sample_rom[130][63] = 8'd130;
	sample_rom[131][0] = 8'd130;
	sample_rom[131][1] = 8'd154;
	sample_rom[131][2] = 8'd172;
	sample_rom[131][3] = 8'd191;
	sample_rom[131][4] = 8'd207;
	sample_rom[131][5] = 8'd222;
	sample_rom[131][6] = 8'd232;
	sample_rom[131][7] = 8'd241;
	sample_rom[131][8] = 8'd246;
	sample_rom[131][9] = 8'd247;
	sample_rom[131][10] = 8'd245;
	sample_rom[131][11] = 8'd240;
	sample_rom[131][12] = 8'd234;
	sample_rom[131][13] = 8'd225;
	sample_rom[131][14] = 8'd215;
	sample_rom[131][15] = 8'd204;
	sample_rom[131][16] = 8'd190;
	sample_rom[131][17] = 8'd176;
	sample_rom[131][18] = 8'd167;
	sample_rom[131][19] = 8'd156;
	sample_rom[131][20] = 8'd145;
	sample_rom[131][21] = 8'd137;
	sample_rom[131][22] = 8'd131;
	sample_rom[131][23] = 8'd127;
	sample_rom[131][24] = 8'd124;
	sample_rom[131][25] = 8'd124;
	sample_rom[131][26] = 8'd123;
	sample_rom[131][27] = 8'd124;
	sample_rom[131][28] = 8'd126;
	sample_rom[131][29] = 8'd130;
	sample_rom[131][30] = 8'd133;
	sample_rom[131][31] = 8'd135;
	sample_rom[131][32] = 8'd138;
	sample_rom[131][33] = 8'd139;
	sample_rom[131][34] = 8'd139;
	sample_rom[131][35] = 8'd138;
	sample_rom[131][36] = 8'd136;
	sample_rom[131][37] = 8'd132;
	sample_rom[131][38] = 8'd129;
	sample_rom[131][39] = 8'd124;
	sample_rom[131][40] = 8'd118;
	sample_rom[131][41] = 8'd114;
	sample_rom[131][42] = 8'd107;
	sample_rom[131][43] = 8'd100;
	sample_rom[131][44] = 8'd96;
	sample_rom[131][45] = 8'd91;
	sample_rom[131][46] = 8'd85;
	sample_rom[131][47] = 8'd81;
	sample_rom[131][48] = 8'd78;
	sample_rom[131][49] = 8'd75;
	sample_rom[131][50] = 8'd76;
	sample_rom[131][51] = 8'd76;
	sample_rom[131][52] = 8'd77;
	sample_rom[131][53] = 8'd80;
	sample_rom[131][54] = 8'd82;
	sample_rom[131][55] = 8'd85;
	sample_rom[131][56] = 8'd90;
	sample_rom[131][57] = 8'd94;
	sample_rom[131][58] = 8'd99;
	sample_rom[131][59] = 8'd104;
	sample_rom[131][60] = 8'd108;
	sample_rom[131][61] = 8'd114;
	sample_rom[131][62] = 8'd119;
	sample_rom[131][63] = 8'd124;
	sample_rom[132][0] = 8'd129;
	sample_rom[132][1] = 8'd187;
	sample_rom[132][2] = 8'd227;
	sample_rom[132][3] = 8'd240;
	sample_rom[132][4] = 8'd230;
	sample_rom[132][5] = 8'd210;
	sample_rom[132][6] = 8'd185;
	sample_rom[132][7] = 8'd173;
	sample_rom[132][8] = 8'd167;
	sample_rom[132][9] = 8'd173;
	sample_rom[132][10] = 8'd181;
	sample_rom[132][11] = 8'd179;
	sample_rom[132][12] = 8'd167;
	sample_rom[132][13] = 8'd150;
	sample_rom[132][14] = 8'd126;
	sample_rom[132][15] = 8'd111;
	sample_rom[132][16] = 8'd103;
	sample_rom[132][17] = 8'd108;
	sample_rom[132][18] = 8'd119;
	sample_rom[132][19] = 8'd127;
	sample_rom[132][20] = 8'd134;
	sample_rom[132][21] = 8'd138;
	sample_rom[132][22] = 8'd140;
	sample_rom[132][23] = 8'd147;
	sample_rom[132][24] = 8'd156;
	sample_rom[132][25] = 8'd166;
	sample_rom[132][26] = 8'd177;
	sample_rom[132][27] = 8'd176;
	sample_rom[132][28] = 8'd170;
	sample_rom[132][29] = 8'd160;
	sample_rom[132][30] = 8'd144;
	sample_rom[132][31] = 8'd130;
	sample_rom[132][32] = 8'd117;
	sample_rom[132][33] = 8'd110;
	sample_rom[132][34] = 8'd107;
	sample_rom[132][35] = 8'd102;
	sample_rom[132][36] = 8'd97;
	sample_rom[132][37] = 8'd94;
	sample_rom[132][38] = 8'd93;
	sample_rom[132][39] = 8'd96;
	sample_rom[132][40] = 8'd103;
	sample_rom[132][41] = 8'd116;
	sample_rom[132][42] = 8'd126;
	sample_rom[132][43] = 8'd133;
	sample_rom[132][44] = 8'd137;
	sample_rom[132][45] = 8'd137;
	sample_rom[132][46] = 8'd138;
	sample_rom[132][47] = 8'd138;
	sample_rom[132][48] = 8'd138;
	sample_rom[132][49] = 8'd138;
	sample_rom[132][50] = 8'd137;
	sample_rom[132][51] = 8'd129;
	sample_rom[132][52] = 8'd120;
	sample_rom[132][53] = 8'd104;
	sample_rom[132][54] = 8'd93;
	sample_rom[132][55] = 8'd85;
	sample_rom[132][56] = 8'd82;
	sample_rom[132][57] = 8'd85;
	sample_rom[132][58] = 8'd91;
	sample_rom[132][59] = 8'd97;
	sample_rom[132][60] = 8'd105;
	sample_rom[132][61] = 8'd113;
	sample_rom[132][62] = 8'd117;
	sample_rom[132][63] = 8'd123;
	sample_rom[133][0] = 8'd128;
	sample_rom[133][1] = 8'd199;
	sample_rom[133][2] = 8'd167;
	sample_rom[133][3] = 8'd208;
	sample_rom[133][4] = 8'd128;
	sample_rom[133][5] = 8'd184;
	sample_rom[133][6] = 8'd146;
	sample_rom[133][7] = 8'd152;
	sample_rom[133][8] = 8'd128;
	sample_rom[133][9] = 8'd162;
	sample_rom[133][10] = 8'd100;
	sample_rom[133][11] = 8'd181;
	sample_rom[133][12] = 8'd128;
	sample_rom[133][13] = 8'd116;
	sample_rom[133][14] = 8'd134;
	sample_rom[133][15] = 8'd98;
	sample_rom[133][16] = 8'd128;
	sample_rom[133][17] = 8'd130;
	sample_rom[133][18] = 8'd140;
	sample_rom[133][19] = 8'd126;
	sample_rom[133][20] = 8'd128;
	sample_rom[133][21] = 8'd188;
	sample_rom[133][22] = 8'd131;
	sample_rom[133][23] = 8'd165;
	sample_rom[133][24] = 8'd128;
	sample_rom[133][25] = 8'd132;
	sample_rom[133][26] = 8'd134;
	sample_rom[133][27] = 8'd182;
	sample_rom[133][28] = 8'd128;
	sample_rom[133][29] = 8'd169;
	sample_rom[133][30] = 8'd150;
	sample_rom[133][31] = 8'd164;
	sample_rom[133][32] = 8'd128;
	sample_rom[133][33] = 8'd94;
	sample_rom[133][34] = 8'd150;
	sample_rom[133][35] = 8'd57;
	sample_rom[133][36] = 8'd128;
	sample_rom[133][37] = 8'd124;
	sample_rom[133][38] = 8'd134;
	sample_rom[133][39] = 8'd82;
	sample_rom[133][40] = 8'd128;
	sample_rom[133][41] = 8'd66;
	sample_rom[133][42] = 8'd131;
	sample_rom[133][43] = 8'd87;
	sample_rom[133][44] = 8'd128;
	sample_rom[133][45] = 8'd151;
	sample_rom[133][46] = 8'd140;
	sample_rom[133][47] = 8'd146;
	sample_rom[133][48] = 8'd128;
	sample_rom[133][49] = 8'd115;
	sample_rom[133][50] = 8'd134;
	sample_rom[133][51] = 8'd147;
	sample_rom[133][52] = 8'd128;
	sample_rom[133][53] = 8'd82;
	sample_rom[133][54] = 8'd100;
	sample_rom[133][55] = 8'd68;
	sample_rom[133][56] = 8'd128;
	sample_rom[133][57] = 8'd102;
	sample_rom[133][58] = 8'd146;
	sample_rom[133][59] = 8'd131;
	sample_rom[133][60] = 8'd128;
	sample_rom[133][61] = 8'd94;
	sample_rom[133][62] = 8'd167;
	sample_rom[133][63] = 8'd128;
	sample_rom[134][0] = 8'd129;
	sample_rom[134][1] = 8'd73;
	sample_rom[134][2] = 8'd84;
	sample_rom[134][3] = 8'd236;
	sample_rom[134][4] = 8'd164;
	sample_rom[134][5] = 8'd168;
	sample_rom[134][6] = 8'd163;
	sample_rom[134][7] = 8'd122;
	sample_rom[134][8] = 8'd101;
	sample_rom[134][9] = 8'd128;
	sample_rom[134][10] = 8'd146;
	sample_rom[134][11] = 8'd130;
	sample_rom[134][12] = 8'd123;
	sample_rom[134][13] = 8'd149;
	sample_rom[134][14] = 8'd160;
	sample_rom[134][15] = 8'd127;
	sample_rom[134][16] = 8'd86;
	sample_rom[134][17] = 8'd97;
	sample_rom[134][18] = 8'd126;
	sample_rom[134][19] = 8'd145;
	sample_rom[134][20] = 8'd152;
	sample_rom[134][21] = 8'd168;
	sample_rom[134][22] = 8'd189;
	sample_rom[134][23] = 8'd177;
	sample_rom[134][24] = 8'd147;
	sample_rom[134][25] = 8'd145;
	sample_rom[134][26] = 8'd162;
	sample_rom[134][27] = 8'd156;
	sample_rom[134][28] = 8'd97;
	sample_rom[134][29] = 8'd46;
	sample_rom[134][30] = 8'd53;
	sample_rom[134][31] = 8'd119;
	sample_rom[134][32] = 8'd177;
	sample_rom[134][33] = 8'd180;
	sample_rom[134][34] = 8'd146;
	sample_rom[134][35] = 8'd141;
	sample_rom[134][36] = 8'd182;
	sample_rom[134][37] = 8'd198;
	sample_rom[134][38] = 8'd161;
	sample_rom[134][39] = 8'd106;
	sample_rom[134][40] = 8'd97;
	sample_rom[134][41] = 8'd128;
	sample_rom[134][42] = 8'd154;
	sample_rom[134][43] = 8'd155;
	sample_rom[134][44] = 8'd160;
	sample_rom[134][45] = 8'd170;
	sample_rom[134][46] = 8'd151;
	sample_rom[134][47] = 8'd100;
	sample_rom[134][48] = 8'd83;
	sample_rom[134][49] = 8'd113;
	sample_rom[134][50] = 8'd149;
	sample_rom[134][51] = 8'd151;
	sample_rom[134][52] = 8'd142;
	sample_rom[134][53] = 8'd145;
	sample_rom[134][54] = 8'd160;
	sample_rom[134][55] = 8'd159;
	sample_rom[134][56] = 8'd154;
	sample_rom[134][57] = 8'd166;
	sample_rom[134][58] = 8'd158;
	sample_rom[134][59] = 8'd103;
	sample_rom[134][60] = 8'd44;
	sample_rom[134][61] = 8'd62;
	sample_rom[134][62] = 8'd144;
	sample_rom[134][63] = 8'd176;
	sample_rom[135][0] = 8'd137;
	sample_rom[135][1] = 8'd41;
	sample_rom[135][2] = 8'd66;
	sample_rom[135][3] = 8'd97;
	sample_rom[135][4] = 8'd191;
	sample_rom[135][5] = 8'd194;
	sample_rom[135][6] = 8'd188;
	sample_rom[135][7] = 8'd116;
	sample_rom[135][8] = 8'd81;
	sample_rom[135][9] = 8'd125;
	sample_rom[135][10] = 8'd157;
	sample_rom[135][11] = 8'd130;
	sample_rom[135][12] = 8'd119;
	sample_rom[135][13] = 8'd162;
	sample_rom[135][14] = 8'd180;
	sample_rom[135][15] = 8'd126;
	sample_rom[135][16] = 8'd64;
	sample_rom[135][17] = 8'd72;
	sample_rom[135][18] = 8'd125;
	sample_rom[135][19] = 8'd152;
	sample_rom[135][20] = 8'd163;
	sample_rom[135][21] = 8'd195;
	sample_rom[135][22] = 8'd223;
	sample_rom[135][23] = 8'd200;
	sample_rom[135][24] = 8'd160;
	sample_rom[135][25] = 8'd152;
	sample_rom[135][26] = 8'd180;
	sample_rom[135][27] = 8'd166;
	sample_rom[135][28] = 8'd80;
	sample_rom[135][29] = 8'd196;
	sample_rom[135][30] = 8'd206;
	sample_rom[135][31] = 8'd116;
	sample_rom[135][32] = 8'd209;
	sample_rom[135][33] = 8'd208;
	sample_rom[135][34] = 8'd155;
	sample_rom[135][35] = 8'd151;
	sample_rom[135][36] = 8'd208;
	sample_rom[135][37] = 8'd41;
	sample_rom[135][38] = 8'd183;
	sample_rom[135][39] = 8'd95;
	sample_rom[135][40] = 8'd78;
	sample_rom[135][41] = 8'd128;
	sample_rom[135][42] = 8'd166;
	sample_rom[135][43] = 8'd176;
	sample_rom[135][44] = 8'd183;
	sample_rom[135][45] = 8'd196;
	sample_rom[135][46] = 8'd165;
	sample_rom[135][47] = 8'd94;
	sample_rom[135][48] = 8'd57;
	sample_rom[135][49] = 8'd102;
	sample_rom[135][50] = 8'd159;
	sample_rom[135][51] = 8'd164;
	sample_rom[135][52] = 8'd142;
	sample_rom[135][53] = 8'd152;
	sample_rom[135][54] = 8'd180;
	sample_rom[135][55] = 8'd178;
	sample_rom[135][56] = 8'd176;
	sample_rom[135][57] = 8'd190;
	sample_rom[135][58] = 8'd177;
	sample_rom[135][59] = 8'd86;
	sample_rom[135][60] = 8'd192;
	sample_rom[135][61] = 8'd223;
	sample_rom[135][62] = 8'd154;
	sample_rom[135][63] = 8'd209;
	sample_rom[136][0] = 8'd131;
	sample_rom[136][1] = 8'd142;
	sample_rom[136][2] = 8'd152;
	sample_rom[136][3] = 8'd160;
	sample_rom[136][4] = 8'd170;
	sample_rom[136][5] = 8'd176;
	sample_rom[136][6] = 8'd185;
	sample_rom[136][7] = 8'd193;
	sample_rom[136][8] = 8'd197;
	sample_rom[136][9] = 8'd204;
	sample_rom[136][10] = 8'd208;
	sample_rom[136][11] = 8'd212;
	sample_rom[136][12] = 8'd215;
	sample_rom[136][13] = 8'd219;
	sample_rom[136][14] = 8'd220;
	sample_rom[136][15] = 8'd223;
	sample_rom[136][16] = 8'd224;
	sample_rom[136][17] = 8'd225;
	sample_rom[136][18] = 8'd223;
	sample_rom[136][19] = 8'd225;
	sample_rom[136][20] = 8'd224;
	sample_rom[136][21] = 8'd224;
	sample_rom[136][22] = 8'd223;
	sample_rom[136][23] = 8'd225;
	sample_rom[136][24] = 8'd223;
	sample_rom[136][25] = 8'd223;
	sample_rom[136][26] = 8'd219;
	sample_rom[136][27] = 8'd218;
	sample_rom[136][28] = 8'd216;
	sample_rom[136][29] = 8'd212;
	sample_rom[136][30] = 8'd210;
	sample_rom[136][31] = 8'd207;
	sample_rom[136][32] = 8'd203;
	sample_rom[136][33] = 8'd200;
	sample_rom[136][34] = 8'd197;
	sample_rom[136][35] = 8'd194;
	sample_rom[136][36] = 8'd190;
	sample_rom[136][37] = 8'd188;
	sample_rom[136][38] = 8'd185;
	sample_rom[136][39] = 8'd182;
	sample_rom[136][40] = 8'd181;
	sample_rom[136][41] = 8'd179;
	sample_rom[136][42] = 8'd179;
	sample_rom[136][43] = 8'd176;
	sample_rom[136][44] = 8'd176;
	sample_rom[136][45] = 8'd174;
	sample_rom[136][46] = 8'd176;
	sample_rom[136][47] = 8'd173;
	sample_rom[136][48] = 8'd173;
	sample_rom[136][49] = 8'd170;
	sample_rom[136][50] = 8'd170;
	sample_rom[136][51] = 8'd166;
	sample_rom[136][52] = 8'd164;
	sample_rom[136][53] = 8'd162;
	sample_rom[136][54] = 8'd160;
	sample_rom[136][55] = 8'd157;
	sample_rom[136][56] = 8'd154;
	sample_rom[136][57] = 8'd149;
	sample_rom[136][58] = 8'd147;
	sample_rom[136][59] = 8'd145;
	sample_rom[136][60] = 8'd141;
	sample_rom[136][61] = 8'd138;
	sample_rom[136][62] = 8'd133;
	sample_rom[136][63] = 8'd130;
	sample_rom[137][0] = 8'd131;
	sample_rom[137][1] = 8'd148;
	sample_rom[137][2] = 8'd163;
	sample_rom[137][3] = 8'd178;
	sample_rom[137][4] = 8'd188;
	sample_rom[137][5] = 8'd199;
	sample_rom[137][6] = 8'd206;
	sample_rom[137][7] = 8'd213;
	sample_rom[137][8] = 8'd216;
	sample_rom[137][9] = 8'd217;
	sample_rom[137][10] = 8'd218;
	sample_rom[137][11] = 8'd218;
	sample_rom[137][12] = 8'd219;
	sample_rom[137][13] = 8'd219;
	sample_rom[137][14] = 8'd221;
	sample_rom[137][15] = 8'd220;
	sample_rom[137][16] = 8'd221;
	sample_rom[137][17] = 8'd225;
	sample_rom[137][18] = 8'd224;
	sample_rom[137][19] = 8'd227;
	sample_rom[137][20] = 8'd226;
	sample_rom[137][21] = 8'd228;
	sample_rom[137][22] = 8'd226;
	sample_rom[137][23] = 8'd226;
	sample_rom[137][24] = 8'd223;
	sample_rom[137][25] = 8'd220;
	sample_rom[137][26] = 8'd216;
	sample_rom[137][27] = 8'd208;
	sample_rom[137][28] = 8'd204;
	sample_rom[137][29] = 8'd197;
	sample_rom[137][30] = 8'd193;
	sample_rom[137][31] = 8'd188;
	sample_rom[137][32] = 8'd182;
	sample_rom[137][33] = 8'd178;
	sample_rom[137][34] = 8'd174;
	sample_rom[137][35] = 8'd173;
	sample_rom[137][36] = 8'd170;
	sample_rom[137][37] = 8'd168;
	sample_rom[137][38] = 8'd166;
	sample_rom[137][39] = 8'd164;
	sample_rom[137][40] = 8'd163;
	sample_rom[137][41] = 8'd163;
	sample_rom[137][42] = 8'd163;
	sample_rom[137][43] = 8'd161;
	sample_rom[137][44] = 8'd159;
	sample_rom[137][45] = 8'd158;
	sample_rom[137][46] = 8'd159;
	sample_rom[137][47] = 8'd157;
	sample_rom[137][48] = 8'd157;
	sample_rom[137][49] = 8'd156;
	sample_rom[137][50] = 8'd154;
	sample_rom[137][51] = 8'd152;
	sample_rom[137][52] = 8'd152;
	sample_rom[137][53] = 8'd151;
	sample_rom[137][54] = 8'd150;
	sample_rom[137][55] = 8'd147;
	sample_rom[137][56] = 8'd147;
	sample_rom[137][57] = 8'd144;
	sample_rom[137][58] = 8'd142;
	sample_rom[137][59] = 8'd142;
	sample_rom[137][60] = 8'd139;
	sample_rom[137][61] = 8'd137;
	sample_rom[137][62] = 8'd133;
	sample_rom[137][63] = 8'd131;
	sample_rom[138][0] = 8'd131;
	sample_rom[138][1] = 8'd175;
	sample_rom[138][2] = 8'd209;
	sample_rom[138][3] = 8'd220;
	sample_rom[138][4] = 8'd215;
	sample_rom[138][5] = 8'd207;
	sample_rom[138][6] = 8'd196;
	sample_rom[138][7] = 8'd191;
	sample_rom[138][8] = 8'd195;
	sample_rom[138][9] = 8'd202;
	sample_rom[138][10] = 8'd207;
	sample_rom[138][11] = 8'd211;
	sample_rom[138][12] = 8'd210;
	sample_rom[138][13] = 8'd208;
	sample_rom[138][14] = 8'd207;
	sample_rom[138][15] = 8'd207;
	sample_rom[138][16] = 8'd211;
	sample_rom[138][17] = 8'd217;
	sample_rom[138][18] = 8'd220;
	sample_rom[138][19] = 8'd223;
	sample_rom[138][20] = 8'd218;
	sample_rom[138][21] = 8'd209;
	sample_rom[138][22] = 8'd196;
	sample_rom[138][23] = 8'd192;
	sample_rom[138][24] = 8'd182;
	sample_rom[138][25] = 8'd180;
	sample_rom[138][26] = 8'd173;
	sample_rom[138][27] = 8'd165;
	sample_rom[138][28] = 8'd154;
	sample_rom[138][29] = 8'd139;
	sample_rom[138][30] = 8'd127;
	sample_rom[138][31] = 8'd120;
	sample_rom[138][32] = 8'd119;
	sample_rom[138][33] = 8'd122;
	sample_rom[138][34] = 8'd125;
	sample_rom[138][35] = 8'd125;
	sample_rom[138][36] = 8'd125;
	sample_rom[138][37] = 8'd118;
	sample_rom[138][38] = 8'd116;
	sample_rom[138][39] = 8'd111;
	sample_rom[138][40] = 8'd104;
	sample_rom[138][41] = 8'd101;
	sample_rom[138][42] = 8'd97;
	sample_rom[138][43] = 8'd96;
	sample_rom[138][44] = 8'd97;
	sample_rom[138][45] = 8'd99;
	sample_rom[138][46] = 8'd100;
	sample_rom[138][47] = 8'd100;
	sample_rom[138][48] = 8'd98;
	sample_rom[138][49] = 8'd102;
	sample_rom[138][50] = 8'd107;
	sample_rom[138][51] = 8'd115;
	sample_rom[138][52] = 8'd122;
	sample_rom[138][53] = 8'd130;
	sample_rom[138][54] = 8'd132;
	sample_rom[138][55] = 8'd129;
	sample_rom[138][56] = 8'd126;
	sample_rom[138][57] = 8'd121;
	sample_rom[138][58] = 8'd118;
	sample_rom[138][59] = 8'd117;
	sample_rom[138][60] = 8'd117;
	sample_rom[138][61] = 8'd117;
	sample_rom[138][62] = 8'd118;
	sample_rom[138][63] = 8'd122;
	sample_rom[139][0] = 8'd129;
	sample_rom[139][1] = 8'd178;
	sample_rom[139][2] = 8'd215;
	sample_rom[139][3] = 8'd227;
	sample_rom[139][4] = 8'd221;
	sample_rom[139][5] = 8'd209;
	sample_rom[139][6] = 8'd190;
	sample_rom[139][7] = 8'd177;
	sample_rom[139][8] = 8'd177;
	sample_rom[139][9] = 8'd183;
	sample_rom[139][10] = 8'd185;
	sample_rom[139][11] = 8'd184;
	sample_rom[139][12] = 8'd179;
	sample_rom[139][13] = 8'd168;
	sample_rom[139][14] = 8'd160;
	sample_rom[139][15] = 8'd157;
	sample_rom[139][16] = 8'd157;
	sample_rom[139][17] = 8'd158;
	sample_rom[139][18] = 8'd160;
	sample_rom[139][19] = 8'd161;
	sample_rom[139][20] = 8'd157;
	sample_rom[139][21] = 8'd151;
	sample_rom[139][22] = 8'd147;
	sample_rom[139][23] = 8'd147;
	sample_rom[139][24] = 8'd149;
	sample_rom[139][25] = 8'd155;
	sample_rom[139][26] = 8'd160;
	sample_rom[139][27] = 8'd162;
	sample_rom[139][28] = 8'd161;
	sample_rom[139][29] = 8'd158;
	sample_rom[139][30] = 8'd148;
	sample_rom[139][31] = 8'd136;
	sample_rom[139][32] = 8'd125;
	sample_rom[139][33] = 8'd119;
	sample_rom[139][34] = 8'd117;
	sample_rom[139][35] = 8'd120;
	sample_rom[139][36] = 8'd126;
	sample_rom[139][37] = 8'd130;
	sample_rom[139][38] = 8'd131;
	sample_rom[139][39] = 8'd128;
	sample_rom[139][40] = 8'd124;
	sample_rom[139][41] = 8'd117;
	sample_rom[139][42] = 8'd109;
	sample_rom[139][43] = 8'd107;
	sample_rom[139][44] = 8'd106;
	sample_rom[139][45] = 8'd109;
	sample_rom[139][46] = 8'd112;
	sample_rom[139][47] = 8'd117;
	sample_rom[139][48] = 8'd119;
	sample_rom[139][49] = 8'd120;
	sample_rom[139][50] = 8'd119;
	sample_rom[139][51] = 8'd118;
	sample_rom[139][52] = 8'd114;
	sample_rom[139][53] = 8'd116;
	sample_rom[139][54] = 8'd120;
	sample_rom[139][55] = 8'd128;
	sample_rom[139][56] = 8'd135;
	sample_rom[139][57] = 8'd137;
	sample_rom[139][58] = 8'd138;
	sample_rom[139][59] = 8'd128;
	sample_rom[139][60] = 8'd122;
	sample_rom[139][61] = 8'd115;
	sample_rom[139][62] = 8'd117;
	sample_rom[139][63] = 8'd119;
	sample_rom[140][0] = 8'd130;
	sample_rom[140][1] = 8'd222;
	sample_rom[140][2] = 8'd246;
	sample_rom[140][3] = 8'd219;
	sample_rom[140][4] = 8'd211;
	sample_rom[140][5] = 8'd223;
	sample_rom[140][6] = 8'd220;
	sample_rom[140][7] = 8'd194;
	sample_rom[140][8] = 8'd178;
	sample_rom[140][9] = 8'd182;
	sample_rom[140][10] = 8'd182;
	sample_rom[140][11] = 8'd161;
	sample_rom[140][12] = 8'd150;
	sample_rom[140][13] = 8'd145;
	sample_rom[140][14] = 8'd125;
	sample_rom[140][15] = 8'd91;
	sample_rom[140][16] = 8'd66;
	sample_rom[140][17] = 8'd79;
	sample_rom[140][18] = 8'd108;
	sample_rom[140][19] = 8'd125;
	sample_rom[140][20] = 8'd134;
	sample_rom[140][21] = 8'd136;
	sample_rom[140][22] = 8'd147;
	sample_rom[140][23] = 8'd164;
	sample_rom[140][24] = 8'd180;
	sample_rom[140][25] = 8'd186;
	sample_rom[140][26] = 8'd173;
	sample_rom[140][27] = 8'd167;
	sample_rom[140][28] = 8'd170;
	sample_rom[140][29] = 8'd165;
	sample_rom[140][30] = 8'd147;
	sample_rom[140][31] = 8'd122;
	sample_rom[140][32] = 8'd110;
	sample_rom[140][33] = 8'd111;
	sample_rom[140][34] = 8'd93;
	sample_rom[140][35] = 8'd78;
	sample_rom[140][36] = 8'd71;
	sample_rom[140][37] = 8'd84;
	sample_rom[140][38] = 8'd89;
	sample_rom[140][39] = 8'd86;
	sample_rom[140][40] = 8'd88;
	sample_rom[140][41] = 8'd113;
	sample_rom[140][42] = 8'd132;
	sample_rom[140][43] = 8'd145;
	sample_rom[140][44] = 8'd145;
	sample_rom[140][45] = 8'd142;
	sample_rom[140][46] = 8'd139;
	sample_rom[140][47] = 8'd142;
	sample_rom[140][48] = 8'd146;
	sample_rom[140][49] = 8'd143;
	sample_rom[140][50] = 8'd144;
	sample_rom[140][51] = 8'd139;
	sample_rom[140][52] = 8'd129;
	sample_rom[140][53] = 8'd108;
	sample_rom[140][54] = 8'd87;
	sample_rom[140][55] = 8'd81;
	sample_rom[140][56] = 8'd86;
	sample_rom[140][57] = 8'd79;
	sample_rom[140][58] = 8'd70;
	sample_rom[140][59] = 8'd83;
	sample_rom[140][60] = 8'd107;
	sample_rom[140][61] = 8'd118;
	sample_rom[140][62] = 8'd113;
	sample_rom[140][63] = 8'd112;
	sample_rom[141][0] = 8'd128;
	sample_rom[141][1] = 8'd203;
	sample_rom[141][2] = 8'd194;
	sample_rom[141][3] = 8'd198;
	sample_rom[141][4] = 8'd183;
	sample_rom[141][5] = 8'd153;
	sample_rom[141][6] = 8'd143;
	sample_rom[141][7] = 8'd156;
	sample_rom[141][8] = 8'd162;
	sample_rom[141][9] = 8'd167;
	sample_rom[141][10] = 8'd156;
	sample_rom[141][11] = 8'd142;
	sample_rom[141][12] = 8'd125;
	sample_rom[141][13] = 8'd125;
	sample_rom[141][14] = 8'd129;
	sample_rom[141][15] = 8'd122;
	sample_rom[141][16] = 8'd116;
	sample_rom[141][17] = 8'd116;
	sample_rom[141][18] = 8'd103;
	sample_rom[141][19] = 8'd104;
	sample_rom[141][20] = 8'd122;
	sample_rom[141][21] = 8'd137;
	sample_rom[141][22] = 8'd139;
	sample_rom[141][23] = 8'd154;
	sample_rom[141][24] = 8'd162;
	sample_rom[141][25] = 8'd153;
	sample_rom[141][26] = 8'd142;
	sample_rom[141][27] = 8'd145;
	sample_rom[141][28] = 8'd138;
	sample_rom[141][29] = 8'd136;
	sample_rom[141][30] = 8'd150;
	sample_rom[141][31] = 8'd144;
	sample_rom[141][32] = 8'd128;
	sample_rom[141][33] = 8'd112;
	sample_rom[141][34] = 8'd103;
	sample_rom[141][35] = 8'd101;
	sample_rom[141][36] = 8'd112;
	sample_rom[141][37] = 8'd124;
	sample_rom[141][38] = 8'd115;
	sample_rom[141][39] = 8'd99;
	sample_rom[141][40] = 8'd103;
	sample_rom[141][41] = 8'd94;
	sample_rom[141][42] = 8'd89;
	sample_rom[141][43] = 8'd160;
	sample_rom[141][44] = 8'd174;
	sample_rom[141][45] = 8'd150;
	sample_rom[141][46] = 8'd154;
	sample_rom[141][47] = 8'd135;
	sample_rom[141][48] = 8'd116;
	sample_rom[141][49] = 8'd126;
	sample_rom[141][50] = 8'd141;
	sample_rom[141][51] = 8'd144;
	sample_rom[141][52] = 8'd138;
	sample_rom[141][53] = 8'd121;
	sample_rom[141][54] = 8'd104;
	sample_rom[141][55] = 8'd93;
	sample_rom[141][56] = 8'd103;
	sample_rom[141][57] = 8'd113;
	sample_rom[141][58] = 8'd115;
	sample_rom[141][59] = 8'd118;
	sample_rom[141][60] = 8'd116;
	sample_rom[141][61] = 8'd106;
	sample_rom[141][62] = 8'd110;
	sample_rom[141][63] = 8'd127;
	sample_rom[142][0] = 8'd128;
	sample_rom[142][1] = 8'd207;
	sample_rom[142][2] = 8'd183;
	sample_rom[142][3] = 8'd171;
	sample_rom[142][4] = 8'd174;
	sample_rom[142][5] = 8'd144;
	sample_rom[142][6] = 8'd142;
	sample_rom[142][7] = 8'd137;
	sample_rom[142][8] = 8'd135;
	sample_rom[142][9] = 8'd154;
	sample_rom[142][10] = 8'd157;
	sample_rom[142][11] = 8'd123;
	sample_rom[142][12] = 8'd121;
	sample_rom[142][13] = 8'd137;
	sample_rom[142][14] = 8'd138;
	sample_rom[142][15] = 8'd122;
	sample_rom[142][16] = 8'd128;
	sample_rom[142][17] = 8'd105;
	sample_rom[142][18] = 8'd97;
	sample_rom[142][19] = 8'd138;
	sample_rom[142][20] = 8'd126;
	sample_rom[142][21] = 8'd122;
	sample_rom[142][22] = 8'd155;
	sample_rom[142][23] = 8'd137;
	sample_rom[142][24] = 8'd135;
	sample_rom[142][25] = 8'd114;
	sample_rom[142][26] = 8'd159;
	sample_rom[142][27] = 8'd148;
	sample_rom[142][28] = 8'd147;
	sample_rom[142][29] = 8'd133;
	sample_rom[142][30] = 8'd148;
	sample_rom[142][31] = 8'd152;
	sample_rom[142][32] = 8'd128;
	sample_rom[142][33] = 8'd96;
	sample_rom[142][34] = 8'd119;
	sample_rom[142][35] = 8'd101;
	sample_rom[142][36] = 8'd92;
	sample_rom[142][37] = 8'd145;
	sample_rom[142][38] = 8'd135;
	sample_rom[142][39] = 8'd104;
	sample_rom[142][40] = 8'd135;
	sample_rom[142][41] = 8'd109;
	sample_rom[142][42] = 8'd96;
	sample_rom[142][43] = 8'd152;
	sample_rom[142][44] = 8'd167;
	sample_rom[142][45] = 8'd137;
	sample_rom[142][46] = 8'd132;
	sample_rom[142][47] = 8'd140;
	sample_rom[142][48] = 8'd128;
	sample_rom[142][49] = 8'd114;
	sample_rom[142][50] = 8'd127;
	sample_rom[142][51] = 8'd114;
	sample_rom[142][52] = 8'd160;
	sample_rom[142][53] = 8'd132;
	sample_rom[142][54] = 8'd99;
	sample_rom[142][55] = 8'd121;
	sample_rom[142][56] = 8'd135;
	sample_rom[142][57] = 8'd122;
	sample_rom[142][58] = 8'd119;
	sample_rom[142][59] = 8'd122;
	sample_rom[142][60] = 8'd114;
	sample_rom[142][61] = 8'd119;
	sample_rom[142][62] = 8'd108;
	sample_rom[142][63] = 8'd107;
	sample_rom[143][0] = 8'd128;
	sample_rom[143][1] = 8'd205;
	sample_rom[143][2] = 8'd180;
	sample_rom[143][3] = 8'd160;
	sample_rom[143][4] = 8'd152;
	sample_rom[143][5] = 8'd139;
	sample_rom[143][6] = 8'd141;
	sample_rom[143][7] = 8'd138;
	sample_rom[143][8] = 8'd128;
	sample_rom[143][9] = 8'd141;
	sample_rom[143][10] = 8'd186;
	sample_rom[143][11] = 8'd99;
	sample_rom[143][12] = 8'd146;
	sample_rom[143][13] = 8'd124;
	sample_rom[143][14] = 8'd115;
	sample_rom[143][15] = 8'd124;
	sample_rom[143][16] = 8'd128;
	sample_rom[143][17] = 8'd104;
	sample_rom[143][18] = 8'd101;
	sample_rom[143][19] = 8'd132;
	sample_rom[143][20] = 8'd152;
	sample_rom[143][21] = 8'd105;
	sample_rom[143][22] = 8'd162;
	sample_rom[143][23] = 8'd121;
	sample_rom[143][24] = 8'd128;
	sample_rom[143][25] = 8'd113;
	sample_rom[143][26] = 8'd159;
	sample_rom[143][27] = 8'd147;
	sample_rom[143][28] = 8'd114;
	sample_rom[143][29] = 8'd138;
	sample_rom[143][30] = 8'd158;
	sample_rom[143][31] = 8'd149;
	sample_rom[143][32] = 8'd128;
	sample_rom[143][33] = 8'd109;
	sample_rom[143][34] = 8'd88;
	sample_rom[143][35] = 8'd128;
	sample_rom[143][36] = 8'd114;
	sample_rom[143][37] = 8'd146;
	sample_rom[143][38] = 8'd123;
	sample_rom[143][39] = 8'd110;
	sample_rom[143][40] = 8'd128;
	sample_rom[143][41] = 8'd116;
	sample_rom[143][42] = 8'd78;
	sample_rom[143][43] = 8'd188;
	sample_rom[143][44] = 8'd152;
	sample_rom[143][45] = 8'd145;
	sample_rom[143][46] = 8'd121;
	sample_rom[143][47] = 8'd144;
	sample_rom[143][48] = 8'd128;
	sample_rom[143][49] = 8'd97;
	sample_rom[143][50] = 8'd136;
	sample_rom[143][51] = 8'd106;
	sample_rom[143][52] = 8'd146;
	sample_rom[143][53] = 8'd154;
	sample_rom[143][54] = 8'd98;
	sample_rom[143][55] = 8'd127;
	sample_rom[143][56] = 8'd128;
	sample_rom[143][57] = 8'd125;
	sample_rom[143][58] = 8'd107;
	sample_rom[143][59] = 8'd111;
	sample_rom[143][60] = 8'd152;
	sample_rom[143][61] = 8'd117;
	sample_rom[143][62] = 8'd107;
	sample_rom[143][63] = 8'd97;
	sample_rom[144][0] = 8'd128;
	sample_rom[144][1] = 8'd202;
	sample_rom[144][2] = 8'd169;
	sample_rom[144][3] = 8'd212;
	sample_rom[144][4] = 8'd128;
	sample_rom[144][5] = 8'd183;
	sample_rom[144][6] = 8'd144;
	sample_rom[144][7] = 8'd155;
	sample_rom[144][8] = 8'd128;
	sample_rom[144][9] = 8'd164;
	sample_rom[144][10] = 8'd99;
	sample_rom[144][11] = 8'd179;
	sample_rom[144][12] = 8'd128;
	sample_rom[144][13] = 8'd114;
	sample_rom[144][14] = 8'd135;
	sample_rom[144][15] = 8'd103;
	sample_rom[144][16] = 8'd128;
	sample_rom[144][17] = 8'd130;
	sample_rom[144][18] = 8'd141;
	sample_rom[144][19] = 8'd121;
	sample_rom[144][20] = 8'd128;
	sample_rom[144][21] = 8'd185;
	sample_rom[144][22] = 8'd130;
	sample_rom[144][23] = 8'd168;
	sample_rom[144][24] = 8'd128;
	sample_rom[144][25] = 8'd135;
	sample_rom[144][26] = 8'd136;
	sample_rom[144][27] = 8'd178;
	sample_rom[144][28] = 8'd128;
	sample_rom[144][29] = 8'd170;
	sample_rom[144][30] = 8'd155;
	sample_rom[144][31] = 8'd165;
	sample_rom[144][32] = 8'd128;
	sample_rom[144][33] = 8'd93;
	sample_rom[144][34] = 8'd155;
	sample_rom[144][35] = 8'd55;
	sample_rom[144][36] = 8'd128;
	sample_rom[144][37] = 8'd121;
	sample_rom[144][38] = 8'd136;
	sample_rom[144][39] = 8'd79;
	sample_rom[144][40] = 8'd128;
	sample_rom[144][41] = 8'd67;
	sample_rom[144][42] = 8'd130;
	sample_rom[144][43] = 8'd91;
	sample_rom[144][44] = 8'd128;
	sample_rom[144][45] = 8'd149;
	sample_rom[144][46] = 8'd141;
	sample_rom[144][47] = 8'd142;
	sample_rom[144][48] = 8'd128;
	sample_rom[144][49] = 8'd116;
	sample_rom[144][50] = 8'd135;
	sample_rom[144][51] = 8'd147;
	sample_rom[144][52] = 8'd128;
	sample_rom[144][53] = 8'd86;
	sample_rom[144][54] = 8'd99;
	sample_rom[144][55] = 8'd68;
	sample_rom[144][56] = 8'd128;
	sample_rom[144][57] = 8'd101;
	sample_rom[144][58] = 8'd144;
	sample_rom[144][59] = 8'd131;
	sample_rom[144][60] = 8'd128;
	sample_rom[144][61] = 8'd94;
	sample_rom[144][62] = 8'd169;
	sample_rom[144][63] = 8'd129;
	sample_rom[145][0] = 8'd132;
	sample_rom[145][1] = 8'd144;
	sample_rom[145][2] = 8'd157;
	sample_rom[145][3] = 8'd169;
	sample_rom[145][4] = 8'd180;
	sample_rom[145][5] = 8'd192;
	sample_rom[145][6] = 8'd202;
	sample_rom[145][7] = 8'd211;
	sample_rom[145][8] = 8'd218;
	sample_rom[145][9] = 8'd225;
	sample_rom[145][10] = 8'd231;
	sample_rom[145][11] = 8'd236;
	sample_rom[145][12] = 8'd239;
	sample_rom[145][13] = 8'd242;
	sample_rom[145][14] = 8'd244;
	sample_rom[145][15] = 8'd245;
	sample_rom[145][16] = 8'd244;
	sample_rom[145][17] = 8'd243;
	sample_rom[145][18] = 8'd240;
	sample_rom[145][19] = 8'd237;
	sample_rom[145][20] = 8'd233;
	sample_rom[145][21] = 8'd229;
	sample_rom[145][22] = 8'd223;
	sample_rom[145][23] = 8'd220;
	sample_rom[145][24] = 8'd214;
	sample_rom[145][25] = 8'd209;
	sample_rom[145][26] = 8'd206;
	sample_rom[145][27] = 8'd200;
	sample_rom[145][28] = 8'd195;
	sample_rom[145][29] = 8'd190;
	sample_rom[145][30] = 8'd186;
	sample_rom[145][31] = 8'd181;
	sample_rom[145][32] = 8'd177;
	sample_rom[145][33] = 8'd174;
	sample_rom[145][34] = 8'd170;
	sample_rom[145][35] = 8'd167;
	sample_rom[145][36] = 8'd165;
	sample_rom[145][37] = 8'd162;
	sample_rom[145][38] = 8'd161;
	sample_rom[145][39] = 8'd159;
	sample_rom[145][40] = 8'd157;
	sample_rom[145][41] = 8'd155;
	sample_rom[145][42] = 8'd153;
	sample_rom[145][43] = 8'd153;
	sample_rom[145][44] = 8'd151;
	sample_rom[145][45] = 8'd149;
	sample_rom[145][46] = 8'd148;
	sample_rom[145][47] = 8'd145;
	sample_rom[145][48] = 8'd145;
	sample_rom[145][49] = 8'd144;
	sample_rom[145][50] = 8'd142;
	sample_rom[145][51] = 8'd141;
	sample_rom[145][52] = 8'd139;
	sample_rom[145][53] = 8'd138;
	sample_rom[145][54] = 8'd136;
	sample_rom[145][55] = 8'd135;
	sample_rom[145][56] = 8'd135;
	sample_rom[145][57] = 8'd133;
	sample_rom[145][58] = 8'd133;
	sample_rom[145][59] = 8'd131;
	sample_rom[145][60] = 8'd131;
	sample_rom[145][61] = 8'd130;
	sample_rom[145][62] = 8'd128;
	sample_rom[145][63] = 8'd128;
	sample_rom[146][0] = 8'd131;
	sample_rom[146][1] = 8'd143;
	sample_rom[146][2] = 8'd154;
	sample_rom[146][3] = 8'd164;
	sample_rom[146][4] = 8'd173;
	sample_rom[146][5] = 8'd184;
	sample_rom[146][6] = 8'd192;
	sample_rom[146][7] = 8'd199;
	sample_rom[146][8] = 8'd206;
	sample_rom[146][9] = 8'd211;
	sample_rom[146][10] = 8'd215;
	sample_rom[146][11] = 8'd218;
	sample_rom[146][12] = 8'd221;
	sample_rom[146][13] = 8'd223;
	sample_rom[146][14] = 8'd222;
	sample_rom[146][15] = 8'd222;
	sample_rom[146][16] = 8'd222;
	sample_rom[146][17] = 8'd221;
	sample_rom[146][18] = 8'd219;
	sample_rom[146][19] = 8'd218;
	sample_rom[146][20] = 8'd216;
	sample_rom[146][21] = 8'd214;
	sample_rom[146][22] = 8'd214;
	sample_rom[146][23] = 8'd212;
	sample_rom[146][24] = 8'd210;
	sample_rom[146][25] = 8'd212;
	sample_rom[146][26] = 8'd211;
	sample_rom[146][27] = 8'd213;
	sample_rom[146][28] = 8'd214;
	sample_rom[146][29] = 8'd214;
	sample_rom[146][30] = 8'd217;
	sample_rom[146][31] = 8'd219;
	sample_rom[146][32] = 8'd219;
	sample_rom[146][33] = 8'd221;
	sample_rom[146][34] = 8'd222;
	sample_rom[146][35] = 8'd223;
	sample_rom[146][36] = 8'd223;
	sample_rom[146][37] = 8'd223;
	sample_rom[146][38] = 8'd223;
	sample_rom[146][39] = 8'd221;
	sample_rom[146][40] = 8'd219;
	sample_rom[146][41] = 8'd215;
	sample_rom[146][42] = 8'd212;
	sample_rom[146][43] = 8'd206;
	sample_rom[146][44] = 8'd202;
	sample_rom[146][45] = 8'd195;
	sample_rom[146][46] = 8'd189;
	sample_rom[146][47] = 8'd180;
	sample_rom[146][48] = 8'd175;
	sample_rom[146][49] = 8'd168;
	sample_rom[146][50] = 8'd162;
	sample_rom[146][51] = 8'd156;
	sample_rom[146][52] = 8'd150;
	sample_rom[146][53] = 8'd144;
	sample_rom[146][54] = 8'd140;
	sample_rom[146][55] = 8'd135;
	sample_rom[146][56] = 8'd132;
	sample_rom[146][57] = 8'd130;
	sample_rom[146][58] = 8'd127;
	sample_rom[146][59] = 8'd126;
	sample_rom[146][60] = 8'd125;
	sample_rom[146][61] = 8'd125;
	sample_rom[146][62] = 8'd125;
	sample_rom[146][63] = 8'd126;
	sample_rom[147][0] = 8'd132;
	sample_rom[147][1] = 8'd149;
	sample_rom[147][2] = 8'd166;
	sample_rom[147][3] = 8'd182;
	sample_rom[147][4] = 8'd196;
	sample_rom[147][5] = 8'd210;
	sample_rom[147][6] = 8'd220;
	sample_rom[147][7] = 8'd228;
	sample_rom[147][8] = 8'd235;
	sample_rom[147][9] = 8'd238;
	sample_rom[147][10] = 8'd241;
	sample_rom[147][11] = 8'd241;
	sample_rom[147][12] = 8'd238;
	sample_rom[147][13] = 8'd233;
	sample_rom[147][14] = 8'd228;
	sample_rom[147][15] = 8'd222;
	sample_rom[147][16] = 8'd215;
	sample_rom[147][17] = 8'd205;
	sample_rom[147][18] = 8'd197;
	sample_rom[147][19] = 8'd189;
	sample_rom[147][20] = 8'd181;
	sample_rom[147][21] = 8'd176;
	sample_rom[147][22] = 8'd169;
	sample_rom[147][23] = 8'd164;
	sample_rom[147][24] = 8'd160;
	sample_rom[147][25] = 8'd157;
	sample_rom[147][26] = 8'd155;
	sample_rom[147][27] = 8'd156;
	sample_rom[147][28] = 8'd154;
	sample_rom[147][29] = 8'd154;
	sample_rom[147][30] = 8'd154;
	sample_rom[147][31] = 8'd155;
	sample_rom[147][32] = 8'd156;
	sample_rom[147][33] = 8'd157;
	sample_rom[147][34] = 8'd157;
	sample_rom[147][35] = 8'd158;
	sample_rom[147][36] = 8'd157;
	sample_rom[147][37] = 8'd155;
	sample_rom[147][38] = 8'd155;
	sample_rom[147][39] = 8'd152;
	sample_rom[147][40] = 8'd152;
	sample_rom[147][41] = 8'd149;
	sample_rom[147][42] = 8'd149;
	sample_rom[147][43] = 8'd146;
	sample_rom[147][44] = 8'd144;
	sample_rom[147][45] = 8'd142;
	sample_rom[147][46] = 8'd140;
	sample_rom[147][47] = 8'd137;
	sample_rom[147][48] = 8'd135;
	sample_rom[147][49] = 8'd134;
	sample_rom[147][50] = 8'd131;
	sample_rom[147][51] = 8'd131;
	sample_rom[147][52] = 8'd132;
	sample_rom[147][53] = 8'd131;
	sample_rom[147][54] = 8'd131;
	sample_rom[147][55] = 8'd131;
	sample_rom[147][56] = 8'd130;
	sample_rom[147][57] = 8'd131;
	sample_rom[147][58] = 8'd131;
	sample_rom[147][59] = 8'd130;
	sample_rom[147][60] = 8'd130;
	sample_rom[147][61] = 8'd128;
	sample_rom[147][62] = 8'd127;
	sample_rom[147][63] = 8'd128;
	sample_rom[148][0] = 8'd130;
	sample_rom[148][1] = 8'd150;
	sample_rom[148][2] = 8'd168;
	sample_rom[148][3] = 8'd184;
	sample_rom[148][4] = 8'd199;
	sample_rom[148][5] = 8'd212;
	sample_rom[148][6] = 8'd223;
	sample_rom[148][7] = 8'd230;
	sample_rom[148][8] = 8'd234;
	sample_rom[148][9] = 8'd237;
	sample_rom[148][10] = 8'd237;
	sample_rom[148][11] = 8'd235;
	sample_rom[148][12] = 8'd229;
	sample_rom[148][13] = 8'd223;
	sample_rom[148][14] = 8'd218;
	sample_rom[148][15] = 8'd211;
	sample_rom[148][16] = 8'd203;
	sample_rom[148][17] = 8'd193;
	sample_rom[148][18] = 8'd187;
	sample_rom[148][19] = 8'd180;
	sample_rom[148][20] = 8'd174;
	sample_rom[148][21] = 8'd168;
	sample_rom[148][22] = 8'd163;
	sample_rom[148][23] = 8'd160;
	sample_rom[148][24] = 8'd156;
	sample_rom[148][25] = 8'd152;
	sample_rom[148][26] = 8'd149;
	sample_rom[148][27] = 8'd147;
	sample_rom[148][28] = 8'd144;
	sample_rom[148][29] = 8'd140;
	sample_rom[148][30] = 8'd136;
	sample_rom[148][31] = 8'd131;
	sample_rom[148][32] = 8'd127;
	sample_rom[148][33] = 8'd122;
	sample_rom[148][34] = 8'd117;
	sample_rom[148][35] = 8'd112;
	sample_rom[148][36] = 8'd106;
	sample_rom[148][37] = 8'd100;
	sample_rom[148][38] = 8'd96;
	sample_rom[148][39] = 8'd93;
	sample_rom[148][40] = 8'd90;
	sample_rom[148][41] = 8'd88;
	sample_rom[148][42] = 8'd87;
	sample_rom[148][43] = 8'd86;
	sample_rom[148][44] = 8'd87;
	sample_rom[148][45] = 8'd89;
	sample_rom[148][46] = 8'd91;
	sample_rom[148][47] = 8'd95;
	sample_rom[148][48] = 8'd97;
	sample_rom[148][49] = 8'd102;
	sample_rom[148][50] = 8'd106;
	sample_rom[148][51] = 8'd110;
	sample_rom[148][52] = 8'd115;
	sample_rom[148][53] = 8'd120;
	sample_rom[148][54] = 8'd123;
	sample_rom[148][55] = 8'd126;
	sample_rom[148][56] = 8'd129;
	sample_rom[148][57] = 8'd130;
	sample_rom[148][58] = 8'd132;
	sample_rom[148][59] = 8'd133;
	sample_rom[148][60] = 8'd132;
	sample_rom[148][61] = 8'd133;
	sample_rom[148][62] = 8'd130;
	sample_rom[148][63] = 8'd129;
	sample_rom[149][0] = 8'd131;
	sample_rom[149][1] = 8'd154;
	sample_rom[149][2] = 8'd174;
	sample_rom[149][3] = 8'd193;
	sample_rom[149][4] = 8'd209;
	sample_rom[149][5] = 8'd223;
	sample_rom[149][6] = 8'd234;
	sample_rom[149][7] = 8'd242;
	sample_rom[149][8] = 8'd245;
	sample_rom[149][9] = 8'd248;
	sample_rom[149][10] = 8'd246;
	sample_rom[149][11] = 8'd245;
	sample_rom[149][12] = 8'd238;
	sample_rom[149][13] = 8'd233;
	sample_rom[149][14] = 8'd228;
	sample_rom[149][15] = 8'd223;
	sample_rom[149][16] = 8'd219;
	sample_rom[149][17] = 8'd213;
	sample_rom[149][18] = 8'd211;
	sample_rom[149][19] = 8'd208;
	sample_rom[149][20] = 8'd209;
	sample_rom[149][21] = 8'd209;
	sample_rom[149][22] = 8'd212;
	sample_rom[149][23] = 8'd215;
	sample_rom[149][24] = 8'd217;
	sample_rom[149][25] = 8'd219;
	sample_rom[149][26] = 8'd220;
	sample_rom[149][27] = 8'd221;
	sample_rom[149][28] = 8'd220;
	sample_rom[149][29] = 8'd219;
	sample_rom[149][30] = 8'd215;
	sample_rom[149][31] = 8'd209;
	sample_rom[149][32] = 8'd205;
	sample_rom[149][33] = 8'd197;
	sample_rom[149][34] = 8'd191;
	sample_rom[149][35] = 8'd184;
	sample_rom[149][36] = 8'd178;
	sample_rom[149][37] = 8'd168;
	sample_rom[149][38] = 8'd163;
	sample_rom[149][39] = 8'd159;
	sample_rom[149][40] = 8'd155;
	sample_rom[149][41] = 8'd152;
	sample_rom[149][42] = 8'd149;
	sample_rom[149][43] = 8'd147;
	sample_rom[149][44] = 8'd147;
	sample_rom[149][45] = 8'd147;
	sample_rom[149][46] = 8'd148;
	sample_rom[149][47] = 8'd148;
	sample_rom[149][48] = 8'd149;
	sample_rom[149][49] = 8'd150;
	sample_rom[149][50] = 8'd151;
	sample_rom[149][51] = 8'd151;
	sample_rom[149][52] = 8'd150;
	sample_rom[149][53] = 8'd149;
	sample_rom[149][54] = 8'd148;
	sample_rom[149][55] = 8'd145;
	sample_rom[149][56] = 8'd142;
	sample_rom[149][57] = 8'd141;
	sample_rom[149][58] = 8'd139;
	sample_rom[149][59] = 8'd137;
	sample_rom[149][60] = 8'd134;
	sample_rom[149][61] = 8'd133;
	sample_rom[149][62] = 8'd130;
	sample_rom[149][63] = 8'd129;
	sample_rom[150][0] = 8'd131;
	sample_rom[150][1] = 8'd151;
	sample_rom[150][2] = 8'd168;
	sample_rom[150][3] = 8'd184;
	sample_rom[150][4] = 8'd198;
	sample_rom[150][5] = 8'd208;
	sample_rom[150][6] = 8'd213;
	sample_rom[150][7] = 8'd218;
	sample_rom[150][8] = 8'd216;
	sample_rom[150][9] = 8'd214;
	sample_rom[150][10] = 8'd210;
	sample_rom[150][11] = 8'd203;
	sample_rom[150][12] = 8'd196;
	sample_rom[150][13] = 8'd187;
	sample_rom[150][14] = 8'd181;
	sample_rom[150][15] = 8'd176;
	sample_rom[150][16] = 8'd171;
	sample_rom[150][17] = 8'd169;
	sample_rom[150][18] = 8'd170;
	sample_rom[150][19] = 8'd172;
	sample_rom[150][20] = 8'd176;
	sample_rom[150][21] = 8'd182;
	sample_rom[150][22] = 8'd187;
	sample_rom[150][23] = 8'd193;
	sample_rom[150][24] = 8'd200;
	sample_rom[150][25] = 8'd206;
	sample_rom[150][26] = 8'd210;
	sample_rom[150][27] = 8'd215;
	sample_rom[150][28] = 8'd216;
	sample_rom[150][29] = 8'd219;
	sample_rom[150][30] = 8'd219;
	sample_rom[150][31] = 8'd219;
	sample_rom[150][32] = 8'd219;
	sample_rom[150][33] = 8'd218;
	sample_rom[150][34] = 8'd218;
	sample_rom[150][35] = 8'd219;
	sample_rom[150][36] = 8'd218;
	sample_rom[150][37] = 8'd221;
	sample_rom[150][38] = 8'd222;
	sample_rom[150][39] = 8'd222;
	sample_rom[150][40] = 8'd224;
	sample_rom[150][41] = 8'd224;
	sample_rom[150][42] = 8'd227;
	sample_rom[150][43] = 8'd224;
	sample_rom[150][44] = 8'd223;
	sample_rom[150][45] = 8'd221;
	sample_rom[150][46] = 8'd217;
	sample_rom[150][47] = 8'd211;
	sample_rom[150][48] = 8'd205;
	sample_rom[150][49] = 8'd196;
	sample_rom[150][50] = 8'd188;
	sample_rom[150][51] = 8'd179;
	sample_rom[150][52] = 8'd169;
	sample_rom[150][53] = 8'd160;
	sample_rom[150][54] = 8'd152;
	sample_rom[150][55] = 8'd144;
	sample_rom[150][56] = 8'd137;
	sample_rom[150][57] = 8'd132;
	sample_rom[150][58] = 8'd128;
	sample_rom[150][59] = 8'd125;
	sample_rom[150][60] = 8'd124;
	sample_rom[150][61] = 8'd123;
	sample_rom[150][62] = 8'd124;
	sample_rom[150][63] = 8'd125;
	sample_rom[151][0] = 8'd132;
	sample_rom[151][1] = 8'd162;
	sample_rom[151][2] = 8'd186;
	sample_rom[151][3] = 8'd209;
	sample_rom[151][4] = 8'd225;
	sample_rom[151][5] = 8'd239;
	sample_rom[151][6] = 8'd247;
	sample_rom[151][7] = 8'd249;
	sample_rom[151][8] = 8'd248;
	sample_rom[151][9] = 8'd240;
	sample_rom[151][10] = 8'd234;
	sample_rom[151][11] = 8'd224;
	sample_rom[151][12] = 8'd216;
	sample_rom[151][13] = 8'd206;
	sample_rom[151][14] = 8'd199;
	sample_rom[151][15] = 8'd195;
	sample_rom[151][16] = 8'd189;
	sample_rom[151][17] = 8'd188;
	sample_rom[151][18] = 8'd187;
	sample_rom[151][19] = 8'd188;
	sample_rom[151][20] = 8'd188;
	sample_rom[151][21] = 8'd188;
	sample_rom[151][22] = 8'd187;
	sample_rom[151][23] = 8'd182;
	sample_rom[151][24] = 8'd177;
	sample_rom[151][25] = 8'd172;
	sample_rom[151][26] = 8'd162;
	sample_rom[151][27] = 8'd157;
	sample_rom[151][28] = 8'd149;
	sample_rom[151][29] = 8'd141;
	sample_rom[151][30] = 8'd136;
	sample_rom[151][31] = 8'd131;
	sample_rom[151][32] = 8'd128;
	sample_rom[151][33] = 8'd128;
	sample_rom[151][34] = 8'd127;
	sample_rom[151][35] = 8'd130;
	sample_rom[151][36] = 8'd132;
	sample_rom[151][37] = 8'd135;
	sample_rom[151][38] = 8'd140;
	sample_rom[151][39] = 8'd140;
	sample_rom[151][40] = 8'd144;
	sample_rom[151][41] = 8'd145;
	sample_rom[151][42] = 8'd144;
	sample_rom[151][43] = 8'd143;
	sample_rom[151][44] = 8'd140;
	sample_rom[151][45] = 8'd138;
	sample_rom[151][46] = 8'd134;
	sample_rom[151][47] = 8'd130;
	sample_rom[151][48] = 8'd126;
	sample_rom[151][49] = 8'd125;
	sample_rom[151][50] = 8'd121;
	sample_rom[151][51] = 8'd121;
	sample_rom[151][52] = 8'd120;
	sample_rom[151][53] = 8'd123;
	sample_rom[151][54] = 8'd123;
	sample_rom[151][55] = 8'd124;
	sample_rom[151][56] = 8'd125;
	sample_rom[151][57] = 8'd127;
	sample_rom[151][58] = 8'd128;
	sample_rom[151][59] = 8'd128;
	sample_rom[151][60] = 8'd130;
	sample_rom[151][61] = 8'd128;
	sample_rom[151][62] = 8'd129;
	sample_rom[151][63] = 8'd129;
	sample_rom[152][0] = 8'd130;
	sample_rom[152][1] = 8'd160;
	sample_rom[152][2] = 8'd186;
	sample_rom[152][3] = 8'd208;
	sample_rom[152][4] = 8'd224;
	sample_rom[152][5] = 8'd236;
	sample_rom[152][6] = 8'd242;
	sample_rom[152][7] = 8'd243;
	sample_rom[152][8] = 8'd238;
	sample_rom[152][9] = 8'd231;
	sample_rom[152][10] = 8'd223;
	sample_rom[152][11] = 8'd215;
	sample_rom[152][12] = 8'd206;
	sample_rom[152][13] = 8'd200;
	sample_rom[152][14] = 8'd195;
	sample_rom[152][15] = 8'd195;
	sample_rom[152][16] = 8'd194;
	sample_rom[152][17] = 8'd194;
	sample_rom[152][18] = 8'd196;
	sample_rom[152][19] = 8'd196;
	sample_rom[152][20] = 8'd195;
	sample_rom[152][21] = 8'd192;
	sample_rom[152][22] = 8'd185;
	sample_rom[152][23] = 8'd178;
	sample_rom[152][24] = 8'd168;
	sample_rom[152][25] = 8'd157;
	sample_rom[152][26] = 8'd145;
	sample_rom[152][27] = 8'd136;
	sample_rom[152][28] = 8'd127;
	sample_rom[152][29] = 8'd120;
	sample_rom[152][30] = 8'd115;
	sample_rom[152][31] = 8'd112;
	sample_rom[152][32] = 8'd111;
	sample_rom[152][33] = 8'd112;
	sample_rom[152][34] = 8'd115;
	sample_rom[152][35] = 8'd116;
	sample_rom[152][36] = 8'd117;
	sample_rom[152][37] = 8'd116;
	sample_rom[152][38] = 8'd113;
	sample_rom[152][39] = 8'd109;
	sample_rom[152][40] = 8'd106;
	sample_rom[152][41] = 8'd99;
	sample_rom[152][42] = 8'd94;
	sample_rom[152][43] = 8'd87;
	sample_rom[152][44] = 8'd83;
	sample_rom[152][45] = 8'd80;
	sample_rom[152][46] = 8'd80;
	sample_rom[152][47] = 8'd82;
	sample_rom[152][48] = 8'd85;
	sample_rom[152][49] = 8'd92;
	sample_rom[152][50] = 8'd98;
	sample_rom[152][51] = 8'd105;
	sample_rom[152][52] = 8'd114;
	sample_rom[152][53] = 8'd122;
	sample_rom[152][54] = 8'd128;
	sample_rom[152][55] = 8'd132;
	sample_rom[152][56] = 8'd137;
	sample_rom[152][57] = 8'd138;
	sample_rom[152][58] = 8'd139;
	sample_rom[152][59] = 8'd140;
	sample_rom[152][60] = 8'd138;
	sample_rom[152][61] = 8'd137;
	sample_rom[152][62] = 8'd133;
	sample_rom[152][63] = 8'd130;
	sample_rom[153][0] = 8'd131;
	sample_rom[153][1] = 8'd168;
	sample_rom[153][2] = 8'd197;
	sample_rom[153][3] = 8'd223;
	sample_rom[153][4] = 8'd236;
	sample_rom[153][5] = 8'd243;
	sample_rom[153][6] = 8'd242;
	sample_rom[153][7] = 8'd233;
	sample_rom[153][8] = 8'd223;
	sample_rom[153][9] = 8'd210;
	sample_rom[153][10] = 8'd202;
	sample_rom[153][11] = 8'd197;
	sample_rom[153][12] = 8'd194;
	sample_rom[153][13] = 8'd199;
	sample_rom[153][14] = 8'd202;
	sample_rom[153][15] = 8'd211;
	sample_rom[153][16] = 8'd217;
	sample_rom[153][17] = 8'd220;
	sample_rom[153][18] = 8'd223;
	sample_rom[153][19] = 8'd222;
	sample_rom[153][20] = 8'd217;
	sample_rom[153][21] = 8'd216;
	sample_rom[153][22] = 8'd212;
	sample_rom[153][23] = 8'd208;
	sample_rom[153][24] = 8'd210;
	sample_rom[153][25] = 8'd210;
	sample_rom[153][26] = 8'd216;
	sample_rom[153][27] = 8'd220;
	sample_rom[153][28] = 8'd227;
	sample_rom[153][29] = 8'd231;
	sample_rom[153][30] = 8'd235;
	sample_rom[153][31] = 8'd237;
	sample_rom[153][32] = 8'd236;
	sample_rom[153][33] = 8'd234;
	sample_rom[153][34] = 8'd229;
	sample_rom[153][35] = 8'd223;
	sample_rom[153][36] = 8'd216;
	sample_rom[153][37] = 8'd208;
	sample_rom[153][38] = 8'd202;
	sample_rom[153][39] = 8'd196;
	sample_rom[153][40] = 8'd189;
	sample_rom[153][41] = 8'd184;
	sample_rom[153][42] = 8'd183;
	sample_rom[153][43] = 8'd180;
	sample_rom[153][44] = 8'd178;
	sample_rom[153][45] = 8'd178;
	sample_rom[153][46] = 8'd179;
	sample_rom[153][47] = 8'd179;
	sample_rom[153][48] = 8'd177;
	sample_rom[153][49] = 8'd175;
	sample_rom[153][50] = 8'd172;
	sample_rom[153][51] = 8'd168;
	sample_rom[153][52] = 8'd160;
	sample_rom[153][53] = 8'd153;
	sample_rom[153][54] = 8'd145;
	sample_rom[153][55] = 8'd136;
	sample_rom[153][56] = 8'd132;
	sample_rom[153][57] = 8'd126;
	sample_rom[153][58] = 8'd123;
	sample_rom[153][59] = 8'd119;
	sample_rom[153][60] = 8'd119;
	sample_rom[153][61] = 8'd118;
	sample_rom[153][62] = 8'd121;
	sample_rom[153][63] = 8'd124;
	sample_rom[154][0] = 8'd131;
	sample_rom[154][1] = 8'd167;
	sample_rom[154][2] = 8'd197;
	sample_rom[154][3] = 8'd221;
	sample_rom[154][4] = 8'd233;
	sample_rom[154][5] = 8'd234;
	sample_rom[154][6] = 8'd229;
	sample_rom[154][7] = 8'd218;
	sample_rom[154][8] = 8'd205;
	sample_rom[154][9] = 8'd194;
	sample_rom[154][10] = 8'd187;
	sample_rom[154][11] = 8'd184;
	sample_rom[154][12] = 8'd184;
	sample_rom[154][13] = 8'd191;
	sample_rom[154][14] = 8'd196;
	sample_rom[154][15] = 8'd202;
	sample_rom[154][16] = 8'd205;
	sample_rom[154][17] = 8'd204;
	sample_rom[154][18] = 8'd201;
	sample_rom[154][19] = 8'd198;
	sample_rom[154][20] = 8'd193;
	sample_rom[154][21] = 8'd189;
	sample_rom[154][22] = 8'd188;
	sample_rom[154][23] = 8'd190;
	sample_rom[154][24] = 8'd189;
	sample_rom[154][25] = 8'd195;
	sample_rom[154][26] = 8'd199;
	sample_rom[154][27] = 8'd203;
	sample_rom[154][28] = 8'd206;
	sample_rom[154][29] = 8'd210;
	sample_rom[154][30] = 8'd210;
	sample_rom[154][31] = 8'd207;
	sample_rom[154][32] = 8'd205;
	sample_rom[154][33] = 8'd202;
	sample_rom[154][34] = 8'd200;
	sample_rom[154][35] = 8'd198;
	sample_rom[154][36] = 8'd197;
	sample_rom[154][37] = 8'd199;
	sample_rom[154][38] = 8'd202;
	sample_rom[154][39] = 8'd205;
	sample_rom[154][40] = 8'd211;
	sample_rom[154][41] = 8'd215;
	sample_rom[154][42] = 8'd220;
	sample_rom[154][43] = 8'd220;
	sample_rom[154][44] = 8'd222;
	sample_rom[154][45] = 8'd219;
	sample_rom[154][46] = 8'd213;
	sample_rom[154][47] = 8'd204;
	sample_rom[154][48] = 8'd198;
	sample_rom[154][49] = 8'd187;
	sample_rom[154][50] = 8'd178;
	sample_rom[154][51] = 8'd167;
	sample_rom[154][52] = 8'd159;
	sample_rom[154][53] = 8'd149;
	sample_rom[154][54] = 8'd143;
	sample_rom[154][55] = 8'd136;
	sample_rom[154][56] = 8'd131;
	sample_rom[154][57] = 8'd129;
	sample_rom[154][58] = 8'd123;
	sample_rom[154][59] = 8'd122;
	sample_rom[154][60] = 8'd120;
	sample_rom[154][61] = 8'd120;
	sample_rom[154][62] = 8'd120;
	sample_rom[154][63] = 8'd125;
	sample_rom[155][0] = 8'd131;
	sample_rom[155][1] = 8'd173;
	sample_rom[155][2] = 8'd210;
	sample_rom[155][3] = 8'd234;
	sample_rom[155][4] = 8'd248;
	sample_rom[155][5] = 8'd252;
	sample_rom[155][6] = 8'd247;
	sample_rom[155][7] = 8'd236;
	sample_rom[155][8] = 8'd226;
	sample_rom[155][9] = 8'd215;
	sample_rom[155][10] = 8'd213;
	sample_rom[155][11] = 8'd213;
	sample_rom[155][12] = 8'd215;
	sample_rom[155][13] = 8'd218;
	sample_rom[155][14] = 8'd217;
	sample_rom[155][15] = 8'd216;
	sample_rom[155][16] = 8'd209;
	sample_rom[155][17] = 8'd201;
	sample_rom[155][18] = 8'd188;
	sample_rom[155][19] = 8'd178;
	sample_rom[155][20] = 8'd171;
	sample_rom[155][21] = 8'd169;
	sample_rom[155][22] = 8'd167;
	sample_rom[155][23] = 8'd168;
	sample_rom[155][24] = 8'd170;
	sample_rom[155][25] = 8'd170;
	sample_rom[155][26] = 8'd167;
	sample_rom[155][27] = 8'd159;
	sample_rom[155][28] = 8'd149;
	sample_rom[155][29] = 8'd139;
	sample_rom[155][30] = 8'd130;
	sample_rom[155][31] = 8'd122;
	sample_rom[155][32] = 8'd115;
	sample_rom[155][33] = 8'd113;
	sample_rom[155][34] = 8'd115;
	sample_rom[155][35] = 8'd118;
	sample_rom[155][36] = 8'd121;
	sample_rom[155][37] = 8'd127;
	sample_rom[155][38] = 8'd128;
	sample_rom[155][39] = 8'd130;
	sample_rom[155][40] = 8'd132;
	sample_rom[155][41] = 8'd133;
	sample_rom[155][42] = 8'd133;
	sample_rom[155][43] = 8'd130;
	sample_rom[155][44] = 8'd128;
	sample_rom[155][45] = 8'd124;
	sample_rom[155][46] = 8'd121;
	sample_rom[155][47] = 8'd118;
	sample_rom[155][48] = 8'd115;
	sample_rom[155][49] = 8'd112;
	sample_rom[155][50] = 8'd111;
	sample_rom[155][51] = 8'd112;
	sample_rom[155][52] = 8'd116;
	sample_rom[155][53] = 8'd119;
	sample_rom[155][54] = 8'd124;
	sample_rom[155][55] = 8'd126;
	sample_rom[155][56] = 8'd132;
	sample_rom[155][57] = 8'd132;
	sample_rom[155][58] = 8'd133;
	sample_rom[155][59] = 8'd133;
	sample_rom[155][60] = 8'd131;
	sample_rom[155][61] = 8'd128;
	sample_rom[155][62] = 8'd128;
	sample_rom[155][63] = 8'd130;
	sample_rom[156][0] = 8'd131;
	sample_rom[156][1] = 8'd178;
	sample_rom[156][2] = 8'd213;
	sample_rom[156][3] = 8'd239;
	sample_rom[156][4] = 8'd248;
	sample_rom[156][5] = 8'd245;
	sample_rom[156][6] = 8'd234;
	sample_rom[156][7] = 8'd223;
	sample_rom[156][8] = 8'd214;
	sample_rom[156][9] = 8'd210;
	sample_rom[156][10] = 8'd213;
	sample_rom[156][11] = 8'd219;
	sample_rom[156][12] = 8'd225;
	sample_rom[156][13] = 8'd229;
	sample_rom[156][14] = 8'd229;
	sample_rom[156][15] = 8'd225;
	sample_rom[156][16] = 8'd222;
	sample_rom[156][17] = 8'd216;
	sample_rom[156][18] = 8'd215;
	sample_rom[156][19] = 8'd215;
	sample_rom[156][20] = 8'd218;
	sample_rom[156][21] = 8'd224;
	sample_rom[156][22] = 8'd223;
	sample_rom[156][23] = 8'd221;
	sample_rom[156][24] = 8'd214;
	sample_rom[156][25] = 8'd203;
	sample_rom[156][26] = 8'd191;
	sample_rom[156][27] = 8'd177;
	sample_rom[156][28] = 8'd166;
	sample_rom[156][29] = 8'd160;
	sample_rom[156][30] = 8'd158;
	sample_rom[156][31] = 8'd157;
	sample_rom[156][32] = 8'd157;
	sample_rom[156][33] = 8'd159;
	sample_rom[156][34] = 8'd157;
	sample_rom[156][35] = 8'd156;
	sample_rom[156][36] = 8'd153;
	sample_rom[156][37] = 8'd146;
	sample_rom[156][38] = 8'd141;
	sample_rom[156][39] = 8'd133;
	sample_rom[156][40] = 8'd125;
	sample_rom[156][41] = 8'd117;
	sample_rom[156][42] = 8'd111;
	sample_rom[156][43] = 8'd104;
	sample_rom[156][44] = 8'd99;
	sample_rom[156][45] = 8'd99;
	sample_rom[156][46] = 8'd100;
	sample_rom[156][47] = 8'd103;
	sample_rom[156][48] = 8'd111;
	sample_rom[156][49] = 8'd118;
	sample_rom[156][50] = 8'd127;
	sample_rom[156][51] = 8'd133;
	sample_rom[156][52] = 8'd141;
	sample_rom[156][53] = 8'd146;
	sample_rom[156][54] = 8'd151;
	sample_rom[156][55] = 8'd154;
	sample_rom[156][56] = 8'd157;
	sample_rom[156][57] = 8'd156;
	sample_rom[156][58] = 8'd156;
	sample_rom[156][59] = 8'd153;
	sample_rom[156][60] = 8'd150;
	sample_rom[156][61] = 8'd147;
	sample_rom[156][62] = 8'd141;
	sample_rom[156][63] = 8'd133;
	sample_rom[157][0] = 8'd131;
	sample_rom[157][1] = 8'd179;
	sample_rom[157][2] = 8'd215;
	sample_rom[157][3] = 8'd236;
	sample_rom[157][4] = 8'd240;
	sample_rom[157][5] = 8'd235;
	sample_rom[157][6] = 8'd222;
	sample_rom[157][7] = 8'd210;
	sample_rom[157][8] = 8'd206;
	sample_rom[157][9] = 8'd203;
	sample_rom[157][10] = 8'd207;
	sample_rom[157][11] = 8'd210;
	sample_rom[157][12] = 8'd209;
	sample_rom[157][13] = 8'd207;
	sample_rom[157][14] = 8'd201;
	sample_rom[157][15] = 8'd196;
	sample_rom[157][16] = 8'd196;
	sample_rom[157][17] = 8'd200;
	sample_rom[157][18] = 8'd206;
	sample_rom[157][19] = 8'd213;
	sample_rom[157][20] = 8'd218;
	sample_rom[157][21] = 8'd220;
	sample_rom[157][22] = 8'd215;
	sample_rom[157][23] = 8'd208;
	sample_rom[157][24] = 8'd203;
	sample_rom[157][25] = 8'd202;
	sample_rom[157][26] = 8'd206;
	sample_rom[157][27] = 8'd216;
	sample_rom[157][28] = 8'd226;
	sample_rom[157][29] = 8'd235;
	sample_rom[157][30] = 8'd246;
	sample_rom[157][31] = 8'd250;
	sample_rom[157][32] = 8'd246;
	sample_rom[157][33] = 8'd241;
	sample_rom[157][34] = 8'd236;
	sample_rom[157][35] = 8'd227;
	sample_rom[157][36] = 8'd219;
	sample_rom[157][37] = 8'd209;
	sample_rom[157][38] = 8'd203;
	sample_rom[157][39] = 8'd195;
	sample_rom[157][40] = 8'd190;
	sample_rom[157][41] = 8'd187;
	sample_rom[157][42] = 8'd191;
	sample_rom[157][43] = 8'd191;
	sample_rom[157][44] = 8'd195;
	sample_rom[157][45] = 8'd195;
	sample_rom[157][46] = 8'd195;
	sample_rom[157][47] = 8'd189;
	sample_rom[157][48] = 8'd184;
	sample_rom[157][49] = 8'd179;
	sample_rom[157][50] = 8'd173;
	sample_rom[157][51] = 8'd167;
	sample_rom[157][52] = 8'd160;
	sample_rom[157][53] = 8'd156;
	sample_rom[157][54] = 8'd150;
	sample_rom[157][55] = 8'd142;
	sample_rom[157][56] = 8'd134;
	sample_rom[157][57] = 8'd127;
	sample_rom[157][58] = 8'd118;
	sample_rom[157][59] = 8'd115;
	sample_rom[157][60] = 8'd112;
	sample_rom[157][61] = 8'd113;
	sample_rom[157][62] = 8'd116;
	sample_rom[157][63] = 8'd121;
	sample_rom[158][0] = 8'd131;
	sample_rom[158][1] = 8'd181;
	sample_rom[158][2] = 8'd216;
	sample_rom[158][3] = 8'd236;
	sample_rom[158][4] = 8'd239;
	sample_rom[158][5] = 8'd228;
	sample_rom[158][6] = 8'd217;
	sample_rom[158][7] = 8'd206;
	sample_rom[158][8] = 8'd203;
	sample_rom[158][9] = 8'd204;
	sample_rom[158][10] = 8'd206;
	sample_rom[158][11] = 8'd204;
	sample_rom[158][12] = 8'd197;
	sample_rom[158][13] = 8'd194;
	sample_rom[158][14] = 8'd191;
	sample_rom[158][15] = 8'd192;
	sample_rom[158][16] = 8'd197;
	sample_rom[158][17] = 8'd204;
	sample_rom[158][18] = 8'd209;
	sample_rom[158][19] = 8'd209;
	sample_rom[158][20] = 8'd203;
	sample_rom[158][21] = 8'd194;
	sample_rom[158][22] = 8'd186;
	sample_rom[158][23] = 8'd183;
	sample_rom[158][24] = 8'd181;
	sample_rom[158][25] = 8'd187;
	sample_rom[158][26] = 8'd194;
	sample_rom[158][27] = 8'd199;
	sample_rom[158][28] = 8'd205;
	sample_rom[158][29] = 8'd210;
	sample_rom[158][30] = 8'd211;
	sample_rom[158][31] = 8'd206;
	sample_rom[158][32] = 8'd203;
	sample_rom[158][33] = 8'd197;
	sample_rom[158][34] = 8'd193;
	sample_rom[158][35] = 8'd190;
	sample_rom[158][36] = 8'd190;
	sample_rom[158][37] = 8'd194;
	sample_rom[158][38] = 8'd200;
	sample_rom[158][39] = 8'd207;
	sample_rom[158][40] = 8'd215;
	sample_rom[158][41] = 8'd220;
	sample_rom[158][42] = 8'd223;
	sample_rom[158][43] = 8'd219;
	sample_rom[158][44] = 8'd219;
	sample_rom[158][45] = 8'd215;
	sample_rom[158][46] = 8'd209;
	sample_rom[158][47] = 8'd206;
	sample_rom[158][48] = 8'd202;
	sample_rom[158][49] = 8'd195;
	sample_rom[158][50] = 8'd185;
	sample_rom[158][51] = 8'd175;
	sample_rom[158][52] = 8'd162;
	sample_rom[158][53] = 8'd152;
	sample_rom[158][54] = 8'd144;
	sample_rom[158][55] = 8'd137;
	sample_rom[158][56] = 8'd132;
	sample_rom[158][57] = 8'd130;
	sample_rom[158][58] = 8'd126;
	sample_rom[158][59] = 8'd125;
	sample_rom[158][60] = 8'd125;
	sample_rom[158][61] = 8'd123;
	sample_rom[158][62] = 8'd123;
	sample_rom[158][63] = 8'd125;
	sample_rom[159][0] = 8'd130;
	sample_rom[159][1] = 8'd185;
	sample_rom[159][2] = 8'd222;
	sample_rom[159][3] = 8'd238;
	sample_rom[159][4] = 8'd238;
	sample_rom[159][5] = 8'd231;
	sample_rom[159][6] = 8'd224;
	sample_rom[159][7] = 8'd222;
	sample_rom[159][8] = 8'd223;
	sample_rom[159][9] = 8'd223;
	sample_rom[159][10] = 8'd217;
	sample_rom[159][11] = 8'd212;
	sample_rom[159][12] = 8'd204;
	sample_rom[159][13] = 8'd202;
	sample_rom[159][14] = 8'd202;
	sample_rom[159][15] = 8'd203;
	sample_rom[159][16] = 8'd200;
	sample_rom[159][17] = 8'd189;
	sample_rom[159][18] = 8'd179;
	sample_rom[159][19] = 8'd169;
	sample_rom[159][20] = 8'd166;
	sample_rom[159][21] = 8'd163;
	sample_rom[159][22] = 8'd165;
	sample_rom[159][23] = 8'd167;
	sample_rom[159][24] = 8'd167;
	sample_rom[159][25] = 8'd162;
	sample_rom[159][26] = 8'd152;
	sample_rom[159][27] = 8'd138;
	sample_rom[159][28] = 8'd122;
	sample_rom[159][29] = 8'd107;
	sample_rom[159][30] = 8'd99;
	sample_rom[159][31] = 8'd95;
	sample_rom[159][32] = 8'd96;
	sample_rom[159][33] = 8'd103;
	sample_rom[159][34] = 8'd107;
	sample_rom[159][35] = 8'd108;
	sample_rom[159][36] = 8'd109;
	sample_rom[159][37] = 8'd104;
	sample_rom[159][38] = 8'd103;
	sample_rom[159][39] = 8'd101;
	sample_rom[159][40] = 8'd98;
	sample_rom[159][41] = 8'd96;
	sample_rom[159][42] = 8'd89;
	sample_rom[159][43] = 8'd84;
	sample_rom[159][44] = 8'd79;
	sample_rom[159][45] = 8'd76;
	sample_rom[159][46] = 8'd75;
	sample_rom[159][47] = 8'd77;
	sample_rom[159][48] = 8'd80;
	sample_rom[159][49] = 8'd84;
	sample_rom[159][50] = 8'd89;
	sample_rom[159][51] = 8'd97;
	sample_rom[159][52] = 8'd104;
	sample_rom[159][53] = 8'd117;
	sample_rom[159][54] = 8'd125;
	sample_rom[159][55] = 8'd130;
	sample_rom[159][56] = 8'd131;
	sample_rom[159][57] = 8'd132;
	sample_rom[159][58] = 8'd135;
	sample_rom[159][59] = 8'd134;
	sample_rom[159][60] = 8'd131;
	sample_rom[159][61] = 8'd132;
	sample_rom[159][62] = 8'd129;
	sample_rom[159][63] = 8'd128;
	sample_rom[160][0] = 8'd132;
	sample_rom[160][1] = 8'd195;
	sample_rom[160][2] = 8'd230;
	sample_rom[160][3] = 8'd245;
	sample_rom[160][4] = 8'd243;
	sample_rom[160][5] = 8'd235;
	sample_rom[160][6] = 8'd231;
	sample_rom[160][7] = 8'd230;
	sample_rom[160][8] = 8'd231;
	sample_rom[160][9] = 8'd229;
	sample_rom[160][10] = 8'd223;
	sample_rom[160][11] = 8'd223;
	sample_rom[160][12] = 8'd227;
	sample_rom[160][13] = 8'd228;
	sample_rom[160][14] = 8'd230;
	sample_rom[160][15] = 8'd229;
	sample_rom[160][16] = 8'd224;
	sample_rom[160][17] = 8'd219;
	sample_rom[160][18] = 8'd218;
	sample_rom[160][19] = 8'd223;
	sample_rom[160][20] = 8'd228;
	sample_rom[160][21] = 8'd231;
	sample_rom[160][22] = 8'd229;
	sample_rom[160][23] = 8'd228;
	sample_rom[160][24] = 8'd221;
	sample_rom[160][25] = 8'd211;
	sample_rom[160][26] = 8'd198;
	sample_rom[160][27] = 8'd182;
	sample_rom[160][28] = 8'd174;
	sample_rom[160][29] = 8'd176;
	sample_rom[160][30] = 8'd179;
	sample_rom[160][31] = 8'd185;
	sample_rom[160][32] = 8'd187;
	sample_rom[160][33] = 8'd187;
	sample_rom[160][34] = 8'd183;
	sample_rom[160][35] = 8'd173;
	sample_rom[160][36] = 8'd169;
	sample_rom[160][37] = 8'd160;
	sample_rom[160][38] = 8'd154;
	sample_rom[160][39] = 8'd146;
	sample_rom[160][40] = 8'd138;
	sample_rom[160][41] = 8'd128;
	sample_rom[160][42] = 8'd124;
	sample_rom[160][43] = 8'd118;
	sample_rom[160][44] = 8'd118;
	sample_rom[160][45] = 8'd120;
	sample_rom[160][46] = 8'd126;
	sample_rom[160][47] = 8'd136;
	sample_rom[160][48] = 8'd141;
	sample_rom[160][49] = 8'd144;
	sample_rom[160][50] = 8'd143;
	sample_rom[160][51] = 8'd141;
	sample_rom[160][52] = 8'd142;
	sample_rom[160][53] = 8'd147;
	sample_rom[160][54] = 8'd150;
	sample_rom[160][55] = 8'd154;
	sample_rom[160][56] = 8'd153;
	sample_rom[160][57] = 8'd153;
	sample_rom[160][58] = 8'd154;
	sample_rom[160][59] = 8'd153;
	sample_rom[160][60] = 8'd148;
	sample_rom[160][61] = 8'd145;
	sample_rom[160][62] = 8'd138;
	sample_rom[160][63] = 8'd133;
	sample_rom[161][0] = 8'd131;
	sample_rom[161][1] = 8'd189;
	sample_rom[161][2] = 8'd223;
	sample_rom[161][3] = 8'd231;
	sample_rom[161][4] = 8'd225;
	sample_rom[161][5] = 8'd220;
	sample_rom[161][6] = 8'd214;
	sample_rom[161][7] = 8'd215;
	sample_rom[161][8] = 8'd209;
	sample_rom[161][9] = 8'd198;
	sample_rom[161][10] = 8'd195;
	sample_rom[161][11] = 8'd200;
	sample_rom[161][12] = 8'd204;
	sample_rom[161][13] = 8'd203;
	sample_rom[161][14] = 8'd198;
	sample_rom[161][15] = 8'd188;
	sample_rom[161][16] = 8'd186;
	sample_rom[161][17] = 8'd195;
	sample_rom[161][18] = 8'd204;
	sample_rom[161][19] = 8'd212;
	sample_rom[161][20] = 8'd215;
	sample_rom[161][21] = 8'd216;
	sample_rom[161][22] = 8'd209;
	sample_rom[161][23] = 8'd204;
	sample_rom[161][24] = 8'd198;
	sample_rom[161][25] = 8'd198;
	sample_rom[161][26] = 8'd205;
	sample_rom[161][27] = 8'd215;
	sample_rom[161][28] = 8'd228;
	sample_rom[161][29] = 8'd239;
	sample_rom[161][30] = 8'd246;
	sample_rom[161][31] = 8'd247;
	sample_rom[161][32] = 8'd248;
	sample_rom[161][33] = 8'd246;
	sample_rom[161][34] = 8'd242;
	sample_rom[161][35] = 8'd233;
	sample_rom[161][36] = 8'd223;
	sample_rom[161][37] = 8'd212;
	sample_rom[161][38] = 8'd206;
	sample_rom[161][39] = 8'd201;
	sample_rom[161][40] = 8'd200;
	sample_rom[161][41] = 8'd198;
	sample_rom[161][42] = 8'd201;
	sample_rom[161][43] = 8'd199;
	sample_rom[161][44] = 8'd200;
	sample_rom[161][45] = 8'd197;
	sample_rom[161][46] = 8'd195;
	sample_rom[161][47] = 8'd192;
	sample_rom[161][48] = 8'd187;
	sample_rom[161][49] = 8'd184;
	sample_rom[161][50] = 8'd178;
	sample_rom[161][51] = 8'd167;
	sample_rom[161][52] = 8'd158;
	sample_rom[161][53] = 8'd151;
	sample_rom[161][54] = 8'd145;
	sample_rom[161][55] = 8'd139;
	sample_rom[161][56] = 8'd129;
	sample_rom[161][57] = 8'd120;
	sample_rom[161][58] = 8'd114;
	sample_rom[161][59] = 8'd111;
	sample_rom[161][60] = 8'd111;
	sample_rom[161][61] = 8'd113;
	sample_rom[161][62] = 8'd114;
	sample_rom[161][63] = 8'd120;
	sample_rom[162][0] = 8'd133;
	sample_rom[162][1] = 8'd190;
	sample_rom[162][2] = 8'd225;
	sample_rom[162][3] = 8'd235;
	sample_rom[162][4] = 8'd233;
	sample_rom[162][5] = 8'd228;
	sample_rom[162][6] = 8'd223;
	sample_rom[162][7] = 8'd223;
	sample_rom[162][8] = 8'd222;
	sample_rom[162][9] = 8'd216;
	sample_rom[162][10] = 8'd215;
	sample_rom[162][11] = 8'd218;
	sample_rom[162][12] = 8'd218;
	sample_rom[162][13] = 8'd213;
	sample_rom[162][14] = 8'd205;
	sample_rom[162][15] = 8'd199;
	sample_rom[162][16] = 8'd204;
	sample_rom[162][17] = 8'd211;
	sample_rom[162][18] = 8'd213;
	sample_rom[162][19] = 8'd207;
	sample_rom[162][20] = 8'd193;
	sample_rom[162][21] = 8'd181;
	sample_rom[162][22] = 8'd172;
	sample_rom[162][23] = 8'd175;
	sample_rom[162][24] = 8'd178;
	sample_rom[162][25] = 8'd182;
	sample_rom[162][26] = 8'd182;
	sample_rom[162][27] = 8'd185;
	sample_rom[162][28] = 8'd185;
	sample_rom[162][29] = 8'd184;
	sample_rom[162][30] = 8'd181;
	sample_rom[162][31] = 8'd171;
	sample_rom[162][32] = 8'd163;
	sample_rom[162][33] = 8'd157;
	sample_rom[162][34] = 8'd148;
	sample_rom[162][35] = 8'd146;
	sample_rom[162][36] = 8'd149;
	sample_rom[162][37] = 8'd157;
	sample_rom[162][38] = 8'd169;
	sample_rom[162][39] = 8'd179;
	sample_rom[162][40] = 8'd184;
	sample_rom[162][41] = 8'd188;
	sample_rom[162][42] = 8'd187;
	sample_rom[162][43] = 8'd187;
	sample_rom[162][44] = 8'd185;
	sample_rom[162][45] = 8'd184;
	sample_rom[162][46] = 8'd178;
	sample_rom[162][47] = 8'd174;
	sample_rom[162][48] = 8'd169;
	sample_rom[162][49] = 8'd162;
	sample_rom[162][50] = 8'd151;
	sample_rom[162][51] = 8'd140;
	sample_rom[162][52] = 8'd127;
	sample_rom[162][53] = 8'd122;
	sample_rom[162][54] = 8'd124;
	sample_rom[162][55] = 8'd125;
	sample_rom[162][56] = 8'd123;
	sample_rom[162][57] = 8'd123;
	sample_rom[162][58] = 8'd123;
	sample_rom[162][59] = 8'd127;
	sample_rom[162][60] = 8'd128;
	sample_rom[162][61] = 8'd129;
	sample_rom[162][62] = 8'd131;
	sample_rom[162][63] = 8'd130;
	sample_rom[163][0] = 8'd130;
	sample_rom[163][1] = 8'd189;
	sample_rom[163][2] = 8'd225;
	sample_rom[163][3] = 8'd241;
	sample_rom[163][4] = 8'd238;
	sample_rom[163][5] = 8'd230;
	sample_rom[163][6] = 8'd223;
	sample_rom[163][7] = 8'd223;
	sample_rom[163][8] = 8'd222;
	sample_rom[163][9] = 8'd221;
	sample_rom[163][10] = 8'd217;
	sample_rom[163][11] = 8'd217;
	sample_rom[163][12] = 8'd212;
	sample_rom[163][13] = 8'd210;
	sample_rom[163][14] = 8'd208;
	sample_rom[163][15] = 8'd209;
	sample_rom[163][16] = 8'd208;
	sample_rom[163][17] = 8'd200;
	sample_rom[163][18] = 8'd191;
	sample_rom[163][19] = 8'd179;
	sample_rom[163][20] = 8'd177;
	sample_rom[163][21] = 8'd176;
	sample_rom[163][22] = 8'd179;
	sample_rom[163][23] = 8'd181;
	sample_rom[163][24] = 8'd176;
	sample_rom[163][25] = 8'd168;
	sample_rom[163][26] = 8'd157;
	sample_rom[163][27] = 8'd145;
	sample_rom[163][28] = 8'd130;
	sample_rom[163][29] = 8'd116;
	sample_rom[163][30] = 8'd106;
	sample_rom[163][31] = 8'd103;
	sample_rom[163][32] = 8'd107;
	sample_rom[163][33] = 8'd116;
	sample_rom[163][34] = 8'd120;
	sample_rom[163][35] = 8'd119;
	sample_rom[163][36] = 8'd118;
	sample_rom[163][37] = 8'd112;
	sample_rom[163][38] = 8'd112;
	sample_rom[163][39] = 8'd110;
	sample_rom[163][40] = 8'd109;
	sample_rom[163][41] = 8'd101;
	sample_rom[163][42] = 8'd96;
	sample_rom[163][43] = 8'd90;
	sample_rom[163][44] = 8'd86;
	sample_rom[163][45] = 8'd79;
	sample_rom[163][46] = 8'd77;
	sample_rom[163][47] = 8'd79;
	sample_rom[163][48] = 8'd83;
	sample_rom[163][49] = 8'd92;
	sample_rom[163][50] = 8'd98;
	sample_rom[163][51] = 8'd105;
	sample_rom[163][52] = 8'd114;
	sample_rom[163][53] = 8'd127;
	sample_rom[163][54] = 8'd134;
	sample_rom[163][55] = 8'd138;
	sample_rom[163][56] = 8'd137;
	sample_rom[163][57] = 8'd134;
	sample_rom[163][58] = 8'd137;
	sample_rom[163][59] = 8'd140;
	sample_rom[163][60] = 8'd137;
	sample_rom[163][61] = 8'd137;
	sample_rom[163][62] = 8'd131;
	sample_rom[163][63] = 8'd127;
	sample_rom[164][0] = 8'd132;
	sample_rom[164][1] = 8'd192;
	sample_rom[164][2] = 8'd228;
	sample_rom[164][3] = 8'd243;
	sample_rom[164][4] = 8'd242;
	sample_rom[164][5] = 8'd235;
	sample_rom[164][6] = 8'd229;
	sample_rom[164][7] = 8'd227;
	sample_rom[164][8] = 8'd229;
	sample_rom[164][9] = 8'd229;
	sample_rom[164][10] = 8'd223;
	sample_rom[164][11] = 8'd222;
	sample_rom[164][12] = 8'd223;
	sample_rom[164][13] = 8'd223;
	sample_rom[164][14] = 8'd225;
	sample_rom[164][15] = 8'd224;
	sample_rom[164][16] = 8'd221;
	sample_rom[164][17] = 8'd214;
	sample_rom[164][18] = 8'd213;
	sample_rom[164][19] = 8'd218;
	sample_rom[164][20] = 8'd224;
	sample_rom[164][21] = 8'd231;
	sample_rom[164][22] = 8'd232;
	sample_rom[164][23] = 8'd232;
	sample_rom[164][24] = 8'd223;
	sample_rom[164][25] = 8'd215;
	sample_rom[164][26] = 8'd204;
	sample_rom[164][27] = 8'd191;
	sample_rom[164][28] = 8'd181;
	sample_rom[164][29] = 8'd180;
	sample_rom[164][30] = 8'd181;
	sample_rom[164][31] = 8'd185;
	sample_rom[164][32] = 8'd189;
	sample_rom[164][33] = 8'd191;
	sample_rom[164][34] = 8'd185;
	sample_rom[164][35] = 8'd175;
	sample_rom[164][36] = 8'd171;
	sample_rom[164][37] = 8'd160;
	sample_rom[164][38] = 8'd156;
	sample_rom[164][39] = 8'd150;
	sample_rom[164][40] = 8'd141;
	sample_rom[164][41] = 8'd128;
	sample_rom[164][42] = 8'd122;
	sample_rom[164][43] = 8'd117;
	sample_rom[164][44] = 8'd117;
	sample_rom[164][45] = 8'd120;
	sample_rom[164][46] = 8'd125;
	sample_rom[164][47] = 8'd134;
	sample_rom[164][48] = 8'd136;
	sample_rom[164][49] = 8'd141;
	sample_rom[164][50] = 8'd142;
	sample_rom[164][51] = 8'd142;
	sample_rom[164][52] = 8'd142;
	sample_rom[164][53] = 8'd145;
	sample_rom[164][54] = 8'd145;
	sample_rom[164][55] = 8'd150;
	sample_rom[164][56] = 8'd150;
	sample_rom[164][57] = 8'd149;
	sample_rom[164][58] = 8'd148;
	sample_rom[164][59] = 8'd145;
	sample_rom[164][60] = 8'd140;
	sample_rom[164][61] = 8'd140;
	sample_rom[164][62] = 8'd137;
	sample_rom[164][63] = 8'd133;
	sample_rom[165][0] = 8'd131;
	sample_rom[165][1] = 8'd190;
	sample_rom[165][2] = 8'd223;
	sample_rom[165][3] = 8'd231;
	sample_rom[165][4] = 8'd227;
	sample_rom[165][5] = 8'd216;
	sample_rom[165][6] = 8'd210;
	sample_rom[165][7] = 8'd208;
	sample_rom[165][8] = 8'd203;
	sample_rom[165][9] = 8'd194;
	sample_rom[165][10] = 8'd192;
	sample_rom[165][11] = 8'd193;
	sample_rom[165][12] = 8'd194;
	sample_rom[165][13] = 8'd193;
	sample_rom[165][14] = 8'd188;
	sample_rom[165][15] = 8'd180;
	sample_rom[165][16] = 8'd185;
	sample_rom[165][17] = 8'd195;
	sample_rom[165][18] = 8'd203;
	sample_rom[165][19] = 8'd209;
	sample_rom[165][20] = 8'd202;
	sample_rom[165][21] = 8'd193;
	sample_rom[165][22] = 8'd185;
	sample_rom[165][23] = 8'd184;
	sample_rom[165][24] = 8'd183;
	sample_rom[165][25] = 8'd190;
	sample_rom[165][26] = 8'd196;
	sample_rom[165][27] = 8'd202;
	sample_rom[165][28] = 8'd207;
	sample_rom[165][29] = 8'd214;
	sample_rom[165][30] = 8'd216;
	sample_rom[165][31] = 8'd211;
	sample_rom[165][32] = 8'd213;
	sample_rom[165][33] = 8'd210;
	sample_rom[165][34] = 8'd206;
	sample_rom[165][35] = 8'd200;
	sample_rom[165][36] = 8'd197;
	sample_rom[165][37] = 8'd199;
	sample_rom[165][38] = 8'd208;
	sample_rom[165][39] = 8'd215;
	sample_rom[165][40] = 8'd223;
	sample_rom[165][41] = 8'd225;
	sample_rom[165][42] = 8'd230;
	sample_rom[165][43] = 8'd227;
	sample_rom[165][44] = 8'd229;
	sample_rom[165][45] = 8'd226;
	sample_rom[165][46] = 8'd219;
	sample_rom[165][47] = 8'd213;
	sample_rom[165][48] = 8'd205;
	sample_rom[165][49] = 8'd198;
	sample_rom[165][50] = 8'd186;
	sample_rom[165][51] = 8'd174;
	sample_rom[165][52] = 8'd163;
	sample_rom[165][53] = 8'd156;
	sample_rom[165][54] = 8'd150;
	sample_rom[165][55] = 8'd144;
	sample_rom[165][56] = 8'd137;
	sample_rom[165][57] = 8'd134;
	sample_rom[165][58] = 8'd129;
	sample_rom[165][59] = 8'd127;
	sample_rom[165][60] = 8'd125;
	sample_rom[165][61] = 8'd122;
	sample_rom[165][62] = 8'd119;
	sample_rom[165][63] = 8'd122;
	sample_rom[166][0] = 8'd132;
	sample_rom[166][1] = 8'd191;
	sample_rom[166][2] = 8'd228;
	sample_rom[166][3] = 8'd242;
	sample_rom[166][4] = 8'd241;
	sample_rom[166][5] = 8'd238;
	sample_rom[166][6] = 8'd233;
	sample_rom[166][7] = 8'd230;
	sample_rom[166][8] = 8'd230;
	sample_rom[166][9] = 8'd222;
	sample_rom[166][10] = 8'd221;
	sample_rom[166][11] = 8'd221;
	sample_rom[166][12] = 8'd216;
	sample_rom[166][13] = 8'd209;
	sample_rom[166][14] = 8'd204;
	sample_rom[166][15] = 8'd200;
	sample_rom[166][16] = 8'd204;
	sample_rom[166][17] = 8'd211;
	sample_rom[166][18] = 8'd206;
	sample_rom[166][19] = 8'd194;
	sample_rom[166][20] = 8'd179;
	sample_rom[166][21] = 8'd171;
	sample_rom[166][22] = 8'd167;
	sample_rom[166][23] = 8'd177;
	sample_rom[166][24] = 8'd179;
	sample_rom[166][25] = 8'd181;
	sample_rom[166][26] = 8'd179;
	sample_rom[166][27] = 8'd177;
	sample_rom[166][28] = 8'd174;
	sample_rom[166][29] = 8'd168;
	sample_rom[166][30] = 8'd158;
	sample_rom[166][31] = 8'd144;
	sample_rom[166][32] = 8'd136;
	sample_rom[166][33] = 8'd130;
	sample_rom[166][34] = 8'd130;
	sample_rom[166][35] = 8'd134;
	sample_rom[166][36] = 8'd139;
	sample_rom[166][37] = 8'd145;
	sample_rom[166][38] = 8'd153;
	sample_rom[166][39] = 8'd159;
	sample_rom[166][40] = 8'd164;
	sample_rom[166][41] = 8'd160;
	sample_rom[166][42] = 8'd161;
	sample_rom[166][43] = 8'd159;
	sample_rom[166][44] = 8'd156;
	sample_rom[166][45] = 8'd155;
	sample_rom[166][46] = 8'd151;
	sample_rom[166][47] = 8'd145;
	sample_rom[166][48] = 8'd141;
	sample_rom[166][49] = 8'd136;
	sample_rom[166][50] = 8'd126;
	sample_rom[166][51] = 8'd122;
	sample_rom[166][52] = 8'd120;
	sample_rom[166][53] = 8'd121;
	sample_rom[166][54] = 8'd122;
	sample_rom[166][55] = 8'd125;
	sample_rom[166][56] = 8'd123;
	sample_rom[166][57] = 8'd124;
	sample_rom[166][58] = 8'd128;
	sample_rom[166][59] = 8'd133;
	sample_rom[166][60] = 8'd133;
	sample_rom[166][61] = 8'd127;
	sample_rom[166][62] = 8'd127;
	sample_rom[166][63] = 8'd127;
	sample_rom[167][0] = 8'd131;
	sample_rom[167][1] = 8'd190;
	sample_rom[167][2] = 8'd227;
	sample_rom[167][3] = 8'd243;
	sample_rom[167][4] = 8'd241;
	sample_rom[167][5] = 8'd234;
	sample_rom[167][6] = 8'd225;
	sample_rom[167][7] = 8'd223;
	sample_rom[167][8] = 8'd223;
	sample_rom[167][9] = 8'd223;
	sample_rom[167][10] = 8'd219;
	sample_rom[167][11] = 8'd220;
	sample_rom[167][12] = 8'd216;
	sample_rom[167][13] = 8'd215;
	sample_rom[167][14] = 8'd216;
	sample_rom[167][15] = 8'd217;
	sample_rom[167][16] = 8'd217;
	sample_rom[167][17] = 8'd211;
	sample_rom[167][18] = 8'd201;
	sample_rom[167][19] = 8'd189;
	sample_rom[167][20] = 8'd187;
	sample_rom[167][21] = 8'd184;
	sample_rom[167][22] = 8'd187;
	sample_rom[167][23] = 8'd189;
	sample_rom[167][24] = 8'd183;
	sample_rom[167][25] = 8'd176;
	sample_rom[167][26] = 8'd165;
	sample_rom[167][27] = 8'd154;
	sample_rom[167][28] = 8'd140;
	sample_rom[167][29] = 8'd127;
	sample_rom[167][30] = 8'd119;
	sample_rom[167][31] = 8'd117;
	sample_rom[167][32] = 8'd121;
	sample_rom[167][33] = 8'd131;
	sample_rom[167][34] = 8'd132;
	sample_rom[167][35] = 8'd130;
	sample_rom[167][36] = 8'd129;
	sample_rom[167][37] = 8'd122;
	sample_rom[167][38] = 8'd120;
	sample_rom[167][39] = 8'd117;
	sample_rom[167][40] = 8'd114;
	sample_rom[167][41] = 8'd107;
	sample_rom[167][42] = 8'd99;
	sample_rom[167][43] = 8'd96;
	sample_rom[167][44] = 8'd91;
	sample_rom[167][45] = 8'd84;
	sample_rom[167][46] = 8'd82;
	sample_rom[167][47] = 8'd83;
	sample_rom[167][48] = 8'd87;
	sample_rom[167][49] = 8'd97;
	sample_rom[167][50] = 8'd103;
	sample_rom[167][51] = 8'd110;
	sample_rom[167][52] = 8'd117;
	sample_rom[167][53] = 8'd132;
	sample_rom[167][54] = 8'd140;
	sample_rom[167][55] = 8'd145;
	sample_rom[167][56] = 8'd143;
	sample_rom[167][57] = 8'd143;
	sample_rom[167][58] = 8'd147;
	sample_rom[167][59] = 8'd149;
	sample_rom[167][60] = 8'd145;
	sample_rom[167][61] = 8'd143;
	sample_rom[167][62] = 8'd137;
	sample_rom[167][63] = 8'd131;
	sample_rom[168][0] = 8'd131;
	sample_rom[168][1] = 8'd194;
	sample_rom[168][2] = 8'd233;
	sample_rom[168][3] = 8'd247;
	sample_rom[168][4] = 8'd245;
	sample_rom[168][5] = 8'd238;
	sample_rom[168][6] = 8'd231;
	sample_rom[168][7] = 8'd229;
	sample_rom[168][8] = 8'd226;
	sample_rom[168][9] = 8'd224;
	sample_rom[168][10] = 8'd219;
	sample_rom[168][11] = 8'd220;
	sample_rom[168][12] = 8'd223;
	sample_rom[168][13] = 8'd224;
	sample_rom[168][14] = 8'd224;
	sample_rom[168][15] = 8'd221;
	sample_rom[168][16] = 8'd214;
	sample_rom[168][17] = 8'd210;
	sample_rom[168][18] = 8'd213;
	sample_rom[168][19] = 8'd222;
	sample_rom[168][20] = 8'd228;
	sample_rom[168][21] = 8'd231;
	sample_rom[168][22] = 8'd231;
	sample_rom[168][23] = 8'd226;
	sample_rom[168][24] = 8'd220;
	sample_rom[168][25] = 8'd212;
	sample_rom[168][26] = 8'd207;
	sample_rom[168][27] = 8'd203;
	sample_rom[168][28] = 8'd204;
	sample_rom[168][29] = 8'd212;
	sample_rom[168][30] = 8'd219;
	sample_rom[168][31] = 8'd223;
	sample_rom[168][32] = 8'd223;
	sample_rom[168][33] = 8'd220;
	sample_rom[168][34] = 8'd217;
	sample_rom[168][35] = 8'd210;
	sample_rom[168][36] = 8'd208;
	sample_rom[168][37] = 8'd201;
	sample_rom[168][38] = 8'd191;
	sample_rom[168][39] = 8'd179;
	sample_rom[168][40] = 8'd170;
	sample_rom[168][41] = 8'd163;
	sample_rom[168][42] = 8'd160;
	sample_rom[168][43] = 8'd160;
	sample_rom[168][44] = 8'd162;
	sample_rom[168][45] = 8'd161;
	sample_rom[168][46] = 8'd164;
	sample_rom[168][47] = 8'd167;
	sample_rom[168][48] = 8'd169;
	sample_rom[168][49] = 8'd164;
	sample_rom[168][50] = 8'd159;
	sample_rom[168][51] = 8'd154;
	sample_rom[168][52] = 8'd154;
	sample_rom[168][53] = 8'd154;
	sample_rom[168][54] = 8'd152;
	sample_rom[168][55] = 8'd150;
	sample_rom[168][56] = 8'd144;
	sample_rom[168][57] = 8'd140;
	sample_rom[168][58] = 8'd139;
	sample_rom[168][59] = 8'd136;
	sample_rom[168][60] = 8'd131;
	sample_rom[168][61] = 8'd131;
	sample_rom[168][62] = 8'd126;
	sample_rom[168][63] = 8'd126;
	sample_rom[169][0] = 8'd131;
	sample_rom[169][1] = 8'd192;
	sample_rom[169][2] = 8'd225;
	sample_rom[169][3] = 8'd236;
	sample_rom[169][4] = 8'd232;
	sample_rom[169][5] = 8'd223;
	sample_rom[169][6] = 8'd220;
	sample_rom[169][7] = 8'd216;
	sample_rom[169][8] = 8'd210;
	sample_rom[169][9] = 8'd201;
	sample_rom[169][10] = 8'd197;
	sample_rom[169][11] = 8'd199;
	sample_rom[169][12] = 8'd200;
	sample_rom[169][13] = 8'd199;
	sample_rom[169][14] = 8'd193;
	sample_rom[169][15] = 8'd187;
	sample_rom[169][16] = 8'd191;
	sample_rom[169][17] = 8'd201;
	sample_rom[169][18] = 8'd210;
	sample_rom[169][19] = 8'd213;
	sample_rom[169][20] = 8'd205;
	sample_rom[169][21] = 8'd194;
	sample_rom[169][22] = 8'd186;
	sample_rom[169][23] = 8'd185;
	sample_rom[169][24] = 8'd183;
	sample_rom[169][25] = 8'd188;
	sample_rom[169][26] = 8'd194;
	sample_rom[169][27] = 8'd199;
	sample_rom[169][28] = 8'd205;
	sample_rom[169][29] = 8'd210;
	sample_rom[169][30] = 8'd208;
	sample_rom[169][31] = 8'd203;
	sample_rom[169][32] = 8'd201;
	sample_rom[169][33] = 8'd197;
	sample_rom[169][34] = 8'd193;
	sample_rom[169][35] = 8'd188;
	sample_rom[169][36] = 8'd187;
	sample_rom[169][37] = 8'd193;
	sample_rom[169][38] = 8'd201;
	sample_rom[169][39] = 8'd211;
	sample_rom[169][40] = 8'd219;
	sample_rom[169][41] = 8'd221;
	sample_rom[169][42] = 8'd222;
	sample_rom[169][43] = 8'd220;
	sample_rom[169][44] = 8'd221;
	sample_rom[169][45] = 8'd216;
	sample_rom[169][46] = 8'd210;
	sample_rom[169][47] = 8'd206;
	sample_rom[169][48] = 8'd201;
	sample_rom[169][49] = 8'd193;
	sample_rom[169][50] = 8'd183;
	sample_rom[169][51] = 8'd173;
	sample_rom[169][52] = 8'd160;
	sample_rom[169][53] = 8'd151;
	sample_rom[169][54] = 8'd144;
	sample_rom[169][55] = 8'd138;
	sample_rom[169][56] = 8'd133;
	sample_rom[169][57] = 8'd130;
	sample_rom[169][58] = 8'd129;
	sample_rom[169][59] = 8'd129;
	sample_rom[169][60] = 8'd128;
	sample_rom[169][61] = 8'd125;
	sample_rom[169][62] = 8'd123;
	sample_rom[169][63] = 8'd123;
	sample_rom[170][0] = 8'd132;
	sample_rom[170][1] = 8'd193;
	sample_rom[170][2] = 8'd231;
	sample_rom[170][3] = 8'd247;
	sample_rom[170][4] = 8'd246;
	sample_rom[170][5] = 8'd242;
	sample_rom[170][6] = 8'd234;
	sample_rom[170][7] = 8'd231;
	sample_rom[170][8] = 8'd229;
	sample_rom[170][9] = 8'd221;
	sample_rom[170][10] = 8'd221;
	sample_rom[170][11] = 8'd222;
	sample_rom[170][12] = 8'd219;
	sample_rom[170][13] = 8'd212;
	sample_rom[170][14] = 8'd207;
	sample_rom[170][15] = 8'd203;
	sample_rom[170][16] = 8'd208;
	sample_rom[170][17] = 8'd213;
	sample_rom[170][18] = 8'd207;
	sample_rom[170][19] = 8'd194;
	sample_rom[170][20] = 8'd178;
	sample_rom[170][21] = 8'd170;
	sample_rom[170][22] = 8'd167;
	sample_rom[170][23] = 8'd176;
	sample_rom[170][24] = 8'd179;
	sample_rom[170][25] = 8'd179;
	sample_rom[170][26] = 8'd176;
	sample_rom[170][27] = 8'd173;
	sample_rom[170][28] = 8'd170;
	sample_rom[170][29] = 8'd164;
	sample_rom[170][30] = 8'd155;
	sample_rom[170][31] = 8'd143;
	sample_rom[170][32] = 8'd136;
	sample_rom[170][33] = 8'd131;
	sample_rom[170][34] = 8'd131;
	sample_rom[170][35] = 8'd136;
	sample_rom[170][36] = 8'd139;
	sample_rom[170][37] = 8'd143;
	sample_rom[170][38] = 8'd149;
	sample_rom[170][39] = 8'd155;
	sample_rom[170][40] = 8'd160;
	sample_rom[170][41] = 8'd158;
	sample_rom[170][42] = 8'd161;
	sample_rom[170][43] = 8'd160;
	sample_rom[170][44] = 8'd160;
	sample_rom[170][45] = 8'd160;
	sample_rom[170][46] = 8'd156;
	sample_rom[170][47] = 8'd148;
	sample_rom[170][48] = 8'd145;
	sample_rom[170][49] = 8'd137;
	sample_rom[170][50] = 8'd125;
	sample_rom[170][51] = 8'd121;
	sample_rom[170][52] = 8'd118;
	sample_rom[170][53] = 8'd120;
	sample_rom[170][54] = 8'd123;
	sample_rom[170][55] = 8'd126;
	sample_rom[170][56] = 8'd126;
	sample_rom[170][57] = 8'd128;
	sample_rom[170][58] = 8'd131;
	sample_rom[170][59] = 8'd135;
	sample_rom[170][60] = 8'd134;
	sample_rom[170][61] = 8'd128;
	sample_rom[170][62] = 8'd127;
	sample_rom[170][63] = 8'd127;
	sample_rom[171][0] = 8'd131;
	sample_rom[171][1] = 8'd188;
	sample_rom[171][2] = 8'd225;
	sample_rom[171][3] = 8'd240;
	sample_rom[171][4] = 8'd241;
	sample_rom[171][5] = 8'd233;
	sample_rom[171][6] = 8'd227;
	sample_rom[171][7] = 8'd227;
	sample_rom[171][8] = 8'd228;
	sample_rom[171][9] = 8'd226;
	sample_rom[171][10] = 8'd221;
	sample_rom[171][11] = 8'd218;
	sample_rom[171][12] = 8'd218;
	sample_rom[171][13] = 8'd220;
	sample_rom[171][14] = 8'd225;
	sample_rom[171][15] = 8'd223;
	sample_rom[171][16] = 8'd222;
	sample_rom[171][17] = 8'd216;
	sample_rom[171][18] = 8'd214;
	sample_rom[171][19] = 8'd217;
	sample_rom[171][20] = 8'd223;
	sample_rom[171][21] = 8'd230;
	sample_rom[171][22] = 8'd230;
	sample_rom[171][23] = 8'd230;
	sample_rom[171][24] = 8'd222;
	sample_rom[171][25] = 8'd213;
	sample_rom[171][26] = 8'd199;
	sample_rom[171][27] = 8'd183;
	sample_rom[171][28] = 8'd170;
	sample_rom[171][29] = 8'd167;
	sample_rom[171][30] = 8'd167;
	sample_rom[171][31] = 8'd172;
	sample_rom[171][32] = 8'd176;
	sample_rom[171][33] = 8'd178;
	sample_rom[171][34] = 8'd173;
	sample_rom[171][35] = 8'd162;
	sample_rom[171][36] = 8'd157;
	sample_rom[171][37] = 8'd148;
	sample_rom[171][38] = 8'd144;
	sample_rom[171][39] = 8'd136;
	sample_rom[171][40] = 8'd127;
	sample_rom[171][41] = 8'd118;
	sample_rom[171][42] = 8'd112;
	sample_rom[171][43] = 8'd108;
	sample_rom[171][44] = 8'd109;
	sample_rom[171][45] = 8'd113;
	sample_rom[171][46] = 8'd115;
	sample_rom[171][47] = 8'd123;
	sample_rom[171][48] = 8'd125;
	sample_rom[171][49] = 8'd133;
	sample_rom[171][50] = 8'd137;
	sample_rom[171][51] = 8'd139;
	sample_rom[171][52] = 8'd142;
	sample_rom[171][53] = 8'd147;
	sample_rom[171][54] = 8'd150;
	sample_rom[171][55] = 8'd154;
	sample_rom[171][56] = 8'd155;
	sample_rom[171][57] = 8'd154;
	sample_rom[171][58] = 8'd155;
	sample_rom[171][59] = 8'd151;
	sample_rom[171][60] = 8'd148;
	sample_rom[171][61] = 8'd148;
	sample_rom[171][62] = 8'd142;
	sample_rom[171][63] = 8'd136;
	sample_rom[172][0] = 8'd131;
	sample_rom[172][1] = 8'd193;
	sample_rom[172][2] = 8'd227;
	sample_rom[172][3] = 8'd241;
	sample_rom[172][4] = 8'd237;
	sample_rom[172][5] = 8'd230;
	sample_rom[172][6] = 8'd227;
	sample_rom[172][7] = 8'd226;
	sample_rom[172][8] = 8'd222;
	sample_rom[172][9] = 8'd214;
	sample_rom[172][10] = 8'd209;
	sample_rom[172][11] = 8'd211;
	sample_rom[172][12] = 8'd214;
	sample_rom[172][13] = 8'd217;
	sample_rom[172][14] = 8'd213;
	sample_rom[172][15] = 8'd206;
	sample_rom[172][16] = 8'd203;
	sample_rom[172][17] = 8'd205;
	sample_rom[172][18] = 8'd213;
	sample_rom[172][19] = 8'd223;
	sample_rom[172][20] = 8'd226;
	sample_rom[172][21] = 8'd230;
	sample_rom[172][22] = 8'd223;
	sample_rom[172][23] = 8'd215;
	sample_rom[172][24] = 8'd208;
	sample_rom[172][25] = 8'd202;
	sample_rom[172][26] = 8'd203;
	sample_rom[172][27] = 8'd205;
	sample_rom[172][28] = 8'd218;
	sample_rom[172][29] = 8'd227;
	sample_rom[172][30] = 8'd236;
	sample_rom[172][31] = 8'd238;
	sample_rom[172][32] = 8'd234;
	sample_rom[172][33] = 8'd231;
	sample_rom[172][34] = 8'd230;
	sample_rom[172][35] = 8'd223;
	sample_rom[172][36] = 8'd217;
	sample_rom[172][37] = 8'd206;
	sample_rom[172][38] = 8'd197;
	sample_rom[172][39] = 8'd187;
	sample_rom[172][40] = 8'd181;
	sample_rom[172][41] = 8'd177;
	sample_rom[172][42] = 8'd180;
	sample_rom[172][43] = 8'd181;
	sample_rom[172][44] = 8'd184;
	sample_rom[172][45] = 8'd186;
	sample_rom[172][46] = 8'd186;
	sample_rom[172][47] = 8'd184;
	sample_rom[172][48] = 8'd179;
	sample_rom[172][49] = 8'd174;
	sample_rom[172][50] = 8'd170;
	sample_rom[172][51] = 8'd168;
	sample_rom[172][52] = 8'd163;
	sample_rom[172][53] = 8'd158;
	sample_rom[172][54] = 8'd150;
	sample_rom[172][55] = 8'd143;
	sample_rom[172][56] = 8'd140;
	sample_rom[172][57] = 8'd131;
	sample_rom[172][58] = 8'd128;
	sample_rom[172][59] = 8'd121;
	sample_rom[172][60] = 8'd118;
	sample_rom[172][61] = 8'd118;
	sample_rom[172][62] = 8'd121;
	sample_rom[172][63] = 8'd124;
	sample_rom[173][0] = 8'd131;
	sample_rom[173][1] = 8'd192;
	sample_rom[173][2] = 8'd224;
	sample_rom[173][3] = 8'd234;
	sample_rom[173][4] = 8'd230;
	sample_rom[173][5] = 8'd223;
	sample_rom[173][6] = 8'd218;
	sample_rom[173][7] = 8'd215;
	sample_rom[173][8] = 8'd211;
	sample_rom[173][9] = 8'd201;
	sample_rom[173][10] = 8'd200;
	sample_rom[173][11] = 8'd202;
	sample_rom[173][12] = 8'd204;
	sample_rom[173][13] = 8'd201;
	sample_rom[173][14] = 8'd197;
	sample_rom[173][15] = 8'd189;
	sample_rom[173][16] = 8'd193;
	sample_rom[173][17] = 8'd204;
	sample_rom[173][18] = 8'd211;
	sample_rom[173][19] = 8'd213;
	sample_rom[173][20] = 8'd204;
	sample_rom[173][21] = 8'd193;
	sample_rom[173][22] = 8'd183;
	sample_rom[173][23] = 8'd181;
	sample_rom[173][24] = 8'd181;
	sample_rom[173][25] = 8'd184;
	sample_rom[173][26] = 8'd189;
	sample_rom[173][27] = 8'd195;
	sample_rom[173][28] = 8'd199;
	sample_rom[173][29] = 8'd202;
	sample_rom[173][30] = 8'd199;
	sample_rom[173][31] = 8'd194;
	sample_rom[173][32] = 8'd191;
	sample_rom[173][33] = 8'd186;
	sample_rom[173][34] = 8'd181;
	sample_rom[173][35] = 8'd176;
	sample_rom[173][36] = 8'd174;
	sample_rom[173][37] = 8'd181;
	sample_rom[173][38] = 8'd192;
	sample_rom[173][39] = 8'd201;
	sample_rom[173][40] = 8'd211;
	sample_rom[173][41] = 8'd212;
	sample_rom[173][42] = 8'd216;
	sample_rom[173][43] = 8'd216;
	sample_rom[173][44] = 8'd216;
	sample_rom[173][45] = 8'd211;
	sample_rom[173][46] = 8'd206;
	sample_rom[173][47] = 8'd202;
	sample_rom[173][48] = 8'd194;
	sample_rom[173][49] = 8'd188;
	sample_rom[173][50] = 8'd177;
	sample_rom[173][51] = 8'd166;
	sample_rom[173][52] = 8'd154;
	sample_rom[173][53] = 8'd145;
	sample_rom[173][54] = 8'd139;
	sample_rom[173][55] = 8'd132;
	sample_rom[173][56] = 8'd126;
	sample_rom[173][57] = 8'd125;
	sample_rom[173][58] = 8'd127;
	sample_rom[173][59] = 8'd128;
	sample_rom[173][60] = 8'd127;
	sample_rom[173][61] = 8'd124;
	sample_rom[173][62] = 8'd124;
	sample_rom[173][63] = 8'd124;
	sample_rom[174][0] = 8'd130;
	sample_rom[174][1] = 8'd193;
	sample_rom[174][2] = 8'd231;
	sample_rom[174][3] = 8'd245;
	sample_rom[174][4] = 8'd245;
	sample_rom[174][5] = 8'd236;
	sample_rom[174][6] = 8'd233;
	sample_rom[174][7] = 8'd227;
	sample_rom[174][8] = 8'd226;
	sample_rom[174][9] = 8'd219;
	sample_rom[174][10] = 8'd215;
	sample_rom[174][11] = 8'd215;
	sample_rom[174][12] = 8'd208;
	sample_rom[174][13] = 8'd202;
	sample_rom[174][14] = 8'd200;
	sample_rom[174][15] = 8'd198;
	sample_rom[174][16] = 8'd203;
	sample_rom[174][17] = 8'd203;
	sample_rom[174][18] = 8'd193;
	sample_rom[174][19] = 8'd176;
	sample_rom[174][20] = 8'd162;
	sample_rom[174][21] = 8'd156;
	sample_rom[174][22] = 8'd157;
	sample_rom[174][23] = 8'd160;
	sample_rom[174][24] = 8'd159;
	sample_rom[174][25] = 8'd155;
	sample_rom[174][26] = 8'd148;
	sample_rom[174][27] = 8'd142;
	sample_rom[174][28] = 8'd135;
	sample_rom[174][29] = 8'd124;
	sample_rom[174][30] = 8'd113;
	sample_rom[174][31] = 8'd100;
	sample_rom[174][32] = 8'd96;
	sample_rom[174][33] = 8'd98;
	sample_rom[174][34] = 8'd103;
	sample_rom[174][35] = 8'd106;
	sample_rom[174][36] = 8'd107;
	sample_rom[174][37] = 8'd107;
	sample_rom[174][38] = 8'd110;
	sample_rom[174][39] = 8'd112;
	sample_rom[174][40] = 8'd111;
	sample_rom[174][41] = 8'd106;
	sample_rom[174][42] = 8'd104;
	sample_rom[174][43] = 8'd102;
	sample_rom[174][44] = 8'd100;
	sample_rom[174][45] = 8'd100;
	sample_rom[174][46] = 8'd96;
	sample_rom[174][47] = 8'd95;
	sample_rom[174][48] = 8'd93;
	sample_rom[174][49] = 8'd97;
	sample_rom[174][50] = 8'd97;
	sample_rom[174][51] = 8'd99;
	sample_rom[174][52] = 8'd102;
	sample_rom[174][53] = 8'd110;
	sample_rom[174][54] = 8'd116;
	sample_rom[174][55] = 8'd124;
	sample_rom[174][56] = 8'd128;
	sample_rom[174][57] = 8'd127;
	sample_rom[174][58] = 8'd126;
	sample_rom[174][59] = 8'd127;
	sample_rom[174][60] = 8'd126;
	sample_rom[174][61] = 8'd126;
	sample_rom[174][62] = 8'd130;
	sample_rom[174][63] = 8'd130;
	sample_rom[175][0] = 8'd130;
	sample_rom[175][1] = 8'd193;
	sample_rom[175][2] = 8'd231;
	sample_rom[175][3] = 8'd245;
	sample_rom[175][4] = 8'd245;
	sample_rom[175][5] = 8'd236;
	sample_rom[175][6] = 8'd233;
	sample_rom[175][7] = 8'd227;
	sample_rom[175][8] = 8'd226;
	sample_rom[175][9] = 8'd219;
	sample_rom[175][10] = 8'd215;
	sample_rom[175][11] = 8'd215;
	sample_rom[175][12] = 8'd208;
	sample_rom[175][13] = 8'd202;
	sample_rom[175][14] = 8'd200;
	sample_rom[175][15] = 8'd198;
	sample_rom[175][16] = 8'd203;
	sample_rom[175][17] = 8'd203;
	sample_rom[175][18] = 8'd193;
	sample_rom[175][19] = 8'd176;
	sample_rom[175][20] = 8'd162;
	sample_rom[175][21] = 8'd156;
	sample_rom[175][22] = 8'd157;
	sample_rom[175][23] = 8'd160;
	sample_rom[175][24] = 8'd159;
	sample_rom[175][25] = 8'd155;
	sample_rom[175][26] = 8'd148;
	sample_rom[175][27] = 8'd142;
	sample_rom[175][28] = 8'd135;
	sample_rom[175][29] = 8'd124;
	sample_rom[175][30] = 8'd113;
	sample_rom[175][31] = 8'd100;
	sample_rom[175][32] = 8'd96;
	sample_rom[175][33] = 8'd98;
	sample_rom[175][34] = 8'd103;
	sample_rom[175][35] = 8'd106;
	sample_rom[175][36] = 8'd107;
	sample_rom[175][37] = 8'd107;
	sample_rom[175][38] = 8'd110;
	sample_rom[175][39] = 8'd112;
	sample_rom[175][40] = 8'd111;
	sample_rom[175][41] = 8'd106;
	sample_rom[175][42] = 8'd104;
	sample_rom[175][43] = 8'd102;
	sample_rom[175][44] = 8'd100;
	sample_rom[175][45] = 8'd100;
	sample_rom[175][46] = 8'd96;
	sample_rom[175][47] = 8'd95;
	sample_rom[175][48] = 8'd93;
	sample_rom[175][49] = 8'd97;
	sample_rom[175][50] = 8'd97;
	sample_rom[175][51] = 8'd99;
	sample_rom[175][52] = 8'd102;
	sample_rom[175][53] = 8'd110;
	sample_rom[175][54] = 8'd116;
	sample_rom[175][55] = 8'd124;
	sample_rom[175][56] = 8'd128;
	sample_rom[175][57] = 8'd127;
	sample_rom[175][58] = 8'd126;
	sample_rom[175][59] = 8'd127;
	sample_rom[175][60] = 8'd126;
	sample_rom[175][61] = 8'd126;
	sample_rom[175][62] = 8'd130;
	sample_rom[175][63] = 8'd130;
	sample_rom[176][0] = 8'd130;
	sample_rom[176][1] = 8'd193;
	sample_rom[176][2] = 8'd231;
	sample_rom[176][3] = 8'd245;
	sample_rom[176][4] = 8'd245;
	sample_rom[176][5] = 8'd236;
	sample_rom[176][6] = 8'd233;
	sample_rom[176][7] = 8'd227;
	sample_rom[176][8] = 8'd226;
	sample_rom[176][9] = 8'd219;
	sample_rom[176][10] = 8'd215;
	sample_rom[176][11] = 8'd215;
	sample_rom[176][12] = 8'd208;
	sample_rom[176][13] = 8'd202;
	sample_rom[176][14] = 8'd200;
	sample_rom[176][15] = 8'd198;
	sample_rom[176][16] = 8'd203;
	sample_rom[176][17] = 8'd203;
	sample_rom[176][18] = 8'd193;
	sample_rom[176][19] = 8'd176;
	sample_rom[176][20] = 8'd162;
	sample_rom[176][21] = 8'd156;
	sample_rom[176][22] = 8'd157;
	sample_rom[176][23] = 8'd160;
	sample_rom[176][24] = 8'd159;
	sample_rom[176][25] = 8'd155;
	sample_rom[176][26] = 8'd148;
	sample_rom[176][27] = 8'd142;
	sample_rom[176][28] = 8'd135;
	sample_rom[176][29] = 8'd124;
	sample_rom[176][30] = 8'd113;
	sample_rom[176][31] = 8'd100;
	sample_rom[176][32] = 8'd96;
	sample_rom[176][33] = 8'd98;
	sample_rom[176][34] = 8'd103;
	sample_rom[176][35] = 8'd106;
	sample_rom[176][36] = 8'd107;
	sample_rom[176][37] = 8'd107;
	sample_rom[176][38] = 8'd110;
	sample_rom[176][39] = 8'd112;
	sample_rom[176][40] = 8'd111;
	sample_rom[176][41] = 8'd106;
	sample_rom[176][42] = 8'd104;
	sample_rom[176][43] = 8'd102;
	sample_rom[176][44] = 8'd100;
	sample_rom[176][45] = 8'd100;
	sample_rom[176][46] = 8'd96;
	sample_rom[176][47] = 8'd95;
	sample_rom[176][48] = 8'd93;
	sample_rom[176][49] = 8'd97;
	sample_rom[176][50] = 8'd97;
	sample_rom[176][51] = 8'd99;
	sample_rom[176][52] = 8'd102;
	sample_rom[176][53] = 8'd110;
	sample_rom[176][54] = 8'd116;
	sample_rom[176][55] = 8'd124;
	sample_rom[176][56] = 8'd128;
	sample_rom[176][57] = 8'd127;
	sample_rom[176][58] = 8'd126;
	sample_rom[176][59] = 8'd127;
	sample_rom[176][60] = 8'd126;
	sample_rom[176][61] = 8'd126;
	sample_rom[176][62] = 8'd130;
	sample_rom[176][63] = 8'd130;
	sample_rom[177][0] = 8'd132;
	sample_rom[177][1] = 8'd150;
	sample_rom[177][2] = 8'd166;
	sample_rom[177][3] = 8'd182;
	sample_rom[177][4] = 8'd197;
	sample_rom[177][5] = 8'd211;
	sample_rom[177][6] = 8'd223;
	sample_rom[177][7] = 8'd232;
	sample_rom[177][8] = 8'd241;
	sample_rom[177][9] = 8'd248;
	sample_rom[177][10] = 8'd253;
	sample_rom[177][11] = 8'd2;
	sample_rom[177][12] = 8'd2;
	sample_rom[177][13] = 8'd252;
	sample_rom[177][14] = 8'd249;
	sample_rom[177][15] = 8'd245;
	sample_rom[177][16] = 8'd238;
	sample_rom[177][17] = 8'd230;
	sample_rom[177][18] = 8'd223;
	sample_rom[177][19] = 8'd215;
	sample_rom[177][20] = 8'd206;
	sample_rom[177][21] = 8'd198;
	sample_rom[177][22] = 8'd189;
	sample_rom[177][23] = 8'd182;
	sample_rom[177][24] = 8'd173;
	sample_rom[177][25] = 8'd168;
	sample_rom[177][26] = 8'd162;
	sample_rom[177][27] = 8'd159;
	sample_rom[177][28] = 8'd156;
	sample_rom[177][29] = 8'd153;
	sample_rom[177][30] = 8'd153;
	sample_rom[177][31] = 8'd152;
	sample_rom[177][32] = 8'd152;
	sample_rom[177][33] = 8'd153;
	sample_rom[177][34] = 8'd153;
	sample_rom[177][35] = 8'd155;
	sample_rom[177][36] = 8'd156;
	sample_rom[177][37] = 8'd157;
	sample_rom[177][38] = 8'd159;
	sample_rom[177][39] = 8'd158;
	sample_rom[177][40] = 8'd160;
	sample_rom[177][41] = 8'd160;
	sample_rom[177][42] = 8'd160;
	sample_rom[177][43] = 8'd157;
	sample_rom[177][44] = 8'd156;
	sample_rom[177][45] = 8'd153;
	sample_rom[177][46] = 8'd151;
	sample_rom[177][47] = 8'd147;
	sample_rom[177][48] = 8'd143;
	sample_rom[177][49] = 8'd141;
	sample_rom[177][50] = 8'd137;
	sample_rom[177][51] = 8'd133;
	sample_rom[177][52] = 8'd130;
	sample_rom[177][53] = 8'd127;
	sample_rom[177][54] = 8'd124;
	sample_rom[177][55] = 8'd122;
	sample_rom[177][56] = 8'd121;
	sample_rom[177][57] = 8'd120;
	sample_rom[177][58] = 8'd120;
	sample_rom[177][59] = 8'd121;
	sample_rom[177][60] = 8'd121;
	sample_rom[177][61] = 8'd122;
	sample_rom[177][62] = 8'd124;
	sample_rom[177][63] = 8'd126;
	sample_rom[178][0] = 8'd132;
	sample_rom[178][1] = 8'd150;
	sample_rom[178][2] = 8'd164;
	sample_rom[178][3] = 8'd180;
	sample_rom[178][4] = 8'd194;
	sample_rom[178][5] = 8'd209;
	sample_rom[178][6] = 8'd220;
	sample_rom[178][7] = 8'd229;
	sample_rom[178][8] = 8'd237;
	sample_rom[178][9] = 8'd243;
	sample_rom[178][10] = 8'd248;
	sample_rom[178][11] = 8'd250;
	sample_rom[178][12] = 8'd249;
	sample_rom[178][13] = 8'd248;
	sample_rom[178][14] = 8'd244;
	sample_rom[178][15] = 8'd240;
	sample_rom[178][16] = 8'd233;
	sample_rom[178][17] = 8'd225;
	sample_rom[178][18] = 8'd220;
	sample_rom[178][19] = 8'd211;
	sample_rom[178][20] = 8'd203;
	sample_rom[178][21] = 8'd195;
	sample_rom[178][22] = 8'd185;
	sample_rom[178][23] = 8'd180;
	sample_rom[178][24] = 8'd172;
	sample_rom[178][25] = 8'd166;
	sample_rom[178][26] = 8'd160;
	sample_rom[178][27] = 8'd157;
	sample_rom[178][28] = 8'd155;
	sample_rom[178][29] = 8'd152;
	sample_rom[178][30] = 8'd153;
	sample_rom[178][31] = 8'd152;
	sample_rom[178][32] = 8'd152;
	sample_rom[178][33] = 8'd153;
	sample_rom[178][34] = 8'd153;
	sample_rom[178][35] = 8'd156;
	sample_rom[178][36] = 8'd157;
	sample_rom[178][37] = 8'd157;
	sample_rom[178][38] = 8'd160;
	sample_rom[178][39] = 8'd159;
	sample_rom[178][40] = 8'd160;
	sample_rom[178][41] = 8'd159;
	sample_rom[178][42] = 8'd160;
	sample_rom[178][43] = 8'd157;
	sample_rom[178][44] = 8'd157;
	sample_rom[178][45] = 8'd154;
	sample_rom[178][46] = 8'd150;
	sample_rom[178][47] = 8'd146;
	sample_rom[178][48] = 8'd143;
	sample_rom[178][49] = 8'd139;
	sample_rom[178][50] = 8'd135;
	sample_rom[178][51] = 8'd132;
	sample_rom[178][52] = 8'd128;
	sample_rom[178][53] = 8'd126;
	sample_rom[178][54] = 8'd124;
	sample_rom[178][55] = 8'd122;
	sample_rom[178][56] = 8'd119;
	sample_rom[178][57] = 8'd120;
	sample_rom[178][58] = 8'd119;
	sample_rom[178][59] = 8'd120;
	sample_rom[178][60] = 8'd120;
	sample_rom[178][61] = 8'd122;
	sample_rom[178][62] = 8'd124;
	sample_rom[178][63] = 8'd126;
	sample_rom[179][0] = 8'd132;
	sample_rom[179][1] = 8'd153;
	sample_rom[179][2] = 8'd172;
	sample_rom[179][3] = 8'd191;
	sample_rom[179][4] = 8'd209;
	sample_rom[179][5] = 8'd223;
	sample_rom[179][6] = 8'd234;
	sample_rom[179][7] = 8'd243;
	sample_rom[179][8] = 8'd250;
	sample_rom[179][9] = 8'd253;
	sample_rom[179][10] = 8'd2;
	sample_rom[179][11] = 8'd251;
	sample_rom[179][12] = 8'd246;
	sample_rom[179][13] = 8'd240;
	sample_rom[179][14] = 8'd231;
	sample_rom[179][15] = 8'd222;
	sample_rom[179][16] = 8'd214;
	sample_rom[179][17] = 8'd203;
	sample_rom[179][18] = 8'd194;
	sample_rom[179][19] = 8'd185;
	sample_rom[179][20] = 8'd177;
	sample_rom[179][21] = 8'd171;
	sample_rom[179][22] = 8'd166;
	sample_rom[179][23] = 8'd164;
	sample_rom[179][24] = 8'd161;
	sample_rom[179][25] = 8'd161;
	sample_rom[179][26] = 8'd160;
	sample_rom[179][27] = 8'd162;
	sample_rom[179][28] = 8'd163;
	sample_rom[179][29] = 8'd165;
	sample_rom[179][30] = 8'd168;
	sample_rom[179][31] = 8'd169;
	sample_rom[179][32] = 8'd171;
	sample_rom[179][33] = 8'd172;
	sample_rom[179][34] = 8'd170;
	sample_rom[179][35] = 8'd170;
	sample_rom[179][36] = 8'd168;
	sample_rom[179][37] = 8'd163;
	sample_rom[179][38] = 8'd161;
	sample_rom[179][39] = 8'd158;
	sample_rom[179][40] = 8'd154;
	sample_rom[179][41] = 8'd149;
	sample_rom[179][42] = 8'd146;
	sample_rom[179][43] = 8'd141;
	sample_rom[179][44] = 8'd138;
	sample_rom[179][45] = 8'd135;
	sample_rom[179][46] = 8'd133;
	sample_rom[179][47] = 8'd130;
	sample_rom[179][48] = 8'd130;
	sample_rom[179][49] = 8'd130;
	sample_rom[179][50] = 8'd131;
	sample_rom[179][51] = 8'd132;
	sample_rom[179][52] = 8'd133;
	sample_rom[179][53] = 8'd136;
	sample_rom[179][54] = 8'd137;
	sample_rom[179][55] = 8'd139;
	sample_rom[179][56] = 8'd137;
	sample_rom[179][57] = 8'd139;
	sample_rom[179][58] = 8'd139;
	sample_rom[179][59] = 8'd137;
	sample_rom[179][60] = 8'd136;
	sample_rom[179][61] = 8'd135;
	sample_rom[179][62] = 8'd133;
	sample_rom[179][63] = 8'd130;
	sample_rom[180][0] = 8'd132;
	sample_rom[180][1] = 8'd156;
	sample_rom[180][2] = 8'd179;
	sample_rom[180][3] = 8'd199;
	sample_rom[180][4] = 8'd217;
	sample_rom[180][5] = 8'd231;
	sample_rom[180][6] = 8'd240;
	sample_rom[180][7] = 8'd246;
	sample_rom[180][8] = 8'd247;
	sample_rom[180][9] = 8'd245;
	sample_rom[180][10] = 8'd241;
	sample_rom[180][11] = 8'd234;
	sample_rom[180][12] = 8'd223;
	sample_rom[180][13] = 8'd212;
	sample_rom[180][14] = 8'd202;
	sample_rom[180][15] = 8'd191;
	sample_rom[180][16] = 8'd182;
	sample_rom[180][17] = 8'd173;
	sample_rom[180][18] = 8'd167;
	sample_rom[180][19] = 8'd163;
	sample_rom[180][20] = 8'd162;
	sample_rom[180][21] = 8'd162;
	sample_rom[180][22] = 8'd162;
	sample_rom[180][23] = 8'd167;
	sample_rom[180][24] = 8'd168;
	sample_rom[180][25] = 8'd172;
	sample_rom[180][26] = 8'd175;
	sample_rom[180][27] = 8'd178;
	sample_rom[180][28] = 8'd178;
	sample_rom[180][29] = 8'd178;
	sample_rom[180][30] = 8'd177;
	sample_rom[180][31] = 8'd174;
	sample_rom[180][32] = 8'd171;
	sample_rom[180][33] = 8'd166;
	sample_rom[180][34] = 8'd160;
	sample_rom[180][35] = 8'd157;
	sample_rom[180][36] = 8'd153;
	sample_rom[180][37] = 8'd147;
	sample_rom[180][38] = 8'd143;
	sample_rom[180][39] = 8'd141;
	sample_rom[180][40] = 8'd141;
	sample_rom[180][41] = 8'd140;
	sample_rom[180][42] = 8'd141;
	sample_rom[180][43] = 8'd142;
	sample_rom[180][44] = 8'd143;
	sample_rom[180][45] = 8'd146;
	sample_rom[180][46] = 8'd146;
	sample_rom[180][47] = 8'd146;
	sample_rom[180][48] = 8'd145;
	sample_rom[180][49] = 8'd146;
	sample_rom[180][50] = 8'd143;
	sample_rom[180][51] = 8'd141;
	sample_rom[180][52] = 8'd137;
	sample_rom[180][53] = 8'd135;
	sample_rom[180][54] = 8'd131;
	sample_rom[180][55] = 8'd127;
	sample_rom[180][56] = 8'd123;
	sample_rom[180][57] = 8'd122;
	sample_rom[180][58] = 8'd120;
	sample_rom[180][59] = 8'd120;
	sample_rom[180][60] = 8'd120;
	sample_rom[180][61] = 8'd121;
	sample_rom[180][62] = 8'd121;
	sample_rom[180][63] = 8'd124;
	sample_rom[181][0] = 8'd132;
	sample_rom[181][1] = 8'd158;
	sample_rom[181][2] = 8'd180;
	sample_rom[181][3] = 8'd202;
	sample_rom[181][4] = 8'd220;
	sample_rom[181][5] = 8'd234;
	sample_rom[181][6] = 8'd245;
	sample_rom[181][7] = 8'd252;
	sample_rom[181][8] = 8'd253;
	sample_rom[181][9] = 8'd252;
	sample_rom[181][10] = 8'd248;
	sample_rom[181][11] = 8'd241;
	sample_rom[181][12] = 8'd230;
	sample_rom[181][13] = 8'd219;
	sample_rom[181][14] = 8'd208;
	sample_rom[181][15] = 8'd197;
	sample_rom[181][16] = 8'd187;
	sample_rom[181][17] = 8'd179;
	sample_rom[181][18] = 8'd171;
	sample_rom[181][19] = 8'd168;
	sample_rom[181][20] = 8'd166;
	sample_rom[181][21] = 8'd165;
	sample_rom[181][22] = 8'd166;
	sample_rom[181][23] = 8'd169;
	sample_rom[181][24] = 8'd170;
	sample_rom[181][25] = 8'd173;
	sample_rom[181][26] = 8'd176;
	sample_rom[181][27] = 8'd177;
	sample_rom[181][28] = 8'd178;
	sample_rom[181][29] = 8'd177;
	sample_rom[181][30] = 8'd176;
	sample_rom[181][31] = 8'd172;
	sample_rom[181][32] = 8'd169;
	sample_rom[181][33] = 8'd163;
	sample_rom[181][34] = 8'd160;
	sample_rom[181][35] = 8'd154;
	sample_rom[181][36] = 8'd149;
	sample_rom[181][37] = 8'd145;
	sample_rom[181][38] = 8'd142;
	sample_rom[181][39] = 8'd139;
	sample_rom[181][40] = 8'd140;
	sample_rom[181][41] = 8'd139;
	sample_rom[181][42] = 8'd140;
	sample_rom[181][43] = 8'd142;
	sample_rom[181][44] = 8'd144;
	sample_rom[181][45] = 8'd146;
	sample_rom[181][46] = 8'd148;
	sample_rom[181][47] = 8'd147;
	sample_rom[181][48] = 8'd147;
	sample_rom[181][49] = 8'd148;
	sample_rom[181][50] = 8'd146;
	sample_rom[181][51] = 8'd144;
	sample_rom[181][52] = 8'd141;
	sample_rom[181][53] = 8'd138;
	sample_rom[181][54] = 8'd134;
	sample_rom[181][55] = 8'd131;
	sample_rom[181][56] = 8'd126;
	sample_rom[181][57] = 8'd125;
	sample_rom[181][58] = 8'd122;
	sample_rom[181][59] = 8'd121;
	sample_rom[181][60] = 8'd122;
	sample_rom[181][61] = 8'd122;
	sample_rom[181][62] = 8'd122;
	sample_rom[181][63] = 8'd125;
	sample_rom[182][0] = 8'd132;
	sample_rom[182][1] = 8'd161;
	sample_rom[182][2] = 8'd189;
	sample_rom[182][3] = 8'd214;
	sample_rom[182][4] = 8'd232;
	sample_rom[182][5] = 8'd247;
	sample_rom[182][6] = 8'd2;
	sample_rom[182][7] = 8'd6;
	sample_rom[182][8] = 8'd2;
	sample_rom[182][9] = 8'd246;
	sample_rom[182][10] = 8'd237;
	sample_rom[182][11] = 8'd224;
	sample_rom[182][12] = 8'd211;
	sample_rom[182][13] = 8'd198;
	sample_rom[182][14] = 8'd187;
	sample_rom[182][15] = 8'd177;
	sample_rom[182][16] = 8'd170;
	sample_rom[182][17] = 8'd167;
	sample_rom[182][18] = 8'd165;
	sample_rom[182][19] = 8'd165;
	sample_rom[182][20] = 8'd169;
	sample_rom[182][21] = 8'd173;
	sample_rom[182][22] = 8'd176;
	sample_rom[182][23] = 8'd180;
	sample_rom[182][24] = 8'd181;
	sample_rom[182][25] = 8'd181;
	sample_rom[182][26] = 8'd179;
	sample_rom[182][27] = 8'd177;
	sample_rom[182][28] = 8'd171;
	sample_rom[182][29] = 8'd166;
	sample_rom[182][30] = 8'd161;
	sample_rom[182][31] = 8'd156;
	sample_rom[182][32] = 8'd152;
	sample_rom[182][33] = 8'd148;
	sample_rom[182][34] = 8'd145;
	sample_rom[182][35] = 8'd145;
	sample_rom[182][36] = 8'd146;
	sample_rom[182][37] = 8'd146;
	sample_rom[182][38] = 8'd148;
	sample_rom[182][39] = 8'd150;
	sample_rom[182][40] = 8'd154;
	sample_rom[182][41] = 8'd154;
	sample_rom[182][42] = 8'd154;
	sample_rom[182][43] = 8'd153;
	sample_rom[182][44] = 8'd151;
	sample_rom[182][45] = 8'd148;
	sample_rom[182][46] = 8'd144;
	sample_rom[182][47] = 8'd138;
	sample_rom[182][48] = 8'd135;
	sample_rom[182][49] = 8'd132;
	sample_rom[182][50] = 8'd128;
	sample_rom[182][51] = 8'd127;
	sample_rom[182][52] = 8'd124;
	sample_rom[182][53] = 8'd127;
	sample_rom[182][54] = 8'd128;
	sample_rom[182][55] = 8'd129;
	sample_rom[182][56] = 8'd131;
	sample_rom[182][57] = 8'd134;
	sample_rom[182][58] = 8'd135;
	sample_rom[182][59] = 8'd136;
	sample_rom[182][60] = 8'd137;
	sample_rom[182][61] = 8'd134;
	sample_rom[182][62] = 8'd132;
	sample_rom[182][63] = 8'd129;
	sample_rom[183][0] = 8'd132;
	sample_rom[183][1] = 8'd166;
	sample_rom[183][2] = 8'd196;
	sample_rom[183][3] = 8'd223;
	sample_rom[183][4] = 8'd242;
	sample_rom[183][5] = 8'd2;
	sample_rom[183][6] = 8'd5;
	sample_rom[183][7] = 8'd4;
	sample_rom[183][8] = 8'd246;
	sample_rom[183][9] = 8'd233;
	sample_rom[183][10] = 8'd221;
	sample_rom[183][11] = 8'd205;
	sample_rom[183][12] = 8'd191;
	sample_rom[183][13] = 8'd180;
	sample_rom[183][14] = 8'd172;
	sample_rom[183][15] = 8'd170;
	sample_rom[183][16] = 8'd168;
	sample_rom[183][17] = 8'd171;
	sample_rom[183][18] = 8'd175;
	sample_rom[183][19] = 8'd179;
	sample_rom[183][20] = 8'd184;
	sample_rom[183][21] = 8'd188;
	sample_rom[183][22] = 8'd189;
	sample_rom[183][23] = 8'd188;
	sample_rom[183][24] = 8'd182;
	sample_rom[183][25] = 8'd177;
	sample_rom[183][26] = 8'd170;
	sample_rom[183][27] = 8'd164;
	sample_rom[183][28] = 8'd159;
	sample_rom[183][29] = 8'd155;
	sample_rom[183][30] = 8'd153;
	sample_rom[183][31] = 8'd150;
	sample_rom[183][32] = 8'd152;
	sample_rom[183][33] = 8'd154;
	sample_rom[183][34] = 8'd156;
	sample_rom[183][35] = 8'd158;
	sample_rom[183][36] = 8'd160;
	sample_rom[183][37] = 8'd160;
	sample_rom[183][38] = 8'd159;
	sample_rom[183][39] = 8'd155;
	sample_rom[183][40] = 8'd155;
	sample_rom[183][41] = 8'd149;
	sample_rom[183][42] = 8'd146;
	sample_rom[183][43] = 8'd142;
	sample_rom[183][44] = 8'd138;
	sample_rom[183][45] = 8'd138;
	sample_rom[183][46] = 8'd136;
	sample_rom[183][47] = 8'd136;
	sample_rom[183][48] = 8'd137;
	sample_rom[183][49] = 8'd140;
	sample_rom[183][50] = 8'd139;
	sample_rom[183][51] = 8'd141;
	sample_rom[183][52] = 8'd139;
	sample_rom[183][53] = 8'd141;
	sample_rom[183][54] = 8'd138;
	sample_rom[183][55] = 8'd135;
	sample_rom[183][56] = 8'd132;
	sample_rom[183][57] = 8'd127;
	sample_rom[183][58] = 8'd124;
	sample_rom[183][59] = 8'd123;
	sample_rom[183][60] = 8'd123;
	sample_rom[183][61] = 8'd122;
	sample_rom[183][62] = 8'd121;
	sample_rom[183][63] = 8'd125;
	sample_rom[184][0] = 8'd131;
	sample_rom[184][1] = 8'd170;
	sample_rom[184][2] = 8'd204;
	sample_rom[184][3] = 8'd232;
	sample_rom[184][4] = 8'd252;
	sample_rom[184][5] = 8'd10;
	sample_rom[184][6] = 8'd8;
	sample_rom[184][7] = 8'd2;
	sample_rom[184][8] = 8'd239;
	sample_rom[184][9] = 8'd223;
	sample_rom[184][10] = 8'd207;
	sample_rom[184][11] = 8'd190;
	sample_rom[184][12] = 8'd179;
	sample_rom[184][13] = 8'd172;
	sample_rom[184][14] = 8'd169;
	sample_rom[184][15] = 8'd171;
	sample_rom[184][16] = 8'd177;
	sample_rom[184][17] = 8'd181;
	sample_rom[184][18] = 8'd186;
	sample_rom[184][19] = 8'd190;
	sample_rom[184][20] = 8'd191;
	sample_rom[184][21] = 8'd189;
	sample_rom[184][22] = 8'd185;
	sample_rom[184][23] = 8'd179;
	sample_rom[184][24] = 8'd172;
	sample_rom[184][25] = 8'd166;
	sample_rom[184][26] = 8'd160;
	sample_rom[184][27] = 8'd158;
	sample_rom[184][28] = 8'd156;
	sample_rom[184][29] = 8'd157;
	sample_rom[184][30] = 8'd160;
	sample_rom[184][31] = 8'd160;
	sample_rom[184][32] = 8'd160;
	sample_rom[184][33] = 8'd161;
	sample_rom[184][34] = 8'd160;
	sample_rom[184][35] = 8'd157;
	sample_rom[184][36] = 8'd153;
	sample_rom[184][37] = 8'd150;
	sample_rom[184][38] = 8'd145;
	sample_rom[184][39] = 8'd141;
	sample_rom[184][40] = 8'd140;
	sample_rom[184][41] = 8'd137;
	sample_rom[184][42] = 8'd139;
	sample_rom[184][43] = 8'd141;
	sample_rom[184][44] = 8'd143;
	sample_rom[184][45] = 8'd145;
	sample_rom[184][46] = 8'd145;
	sample_rom[184][47] = 8'd145;
	sample_rom[184][48] = 8'd144;
	sample_rom[184][49] = 8'd144;
	sample_rom[184][50] = 8'd138;
	sample_rom[184][51] = 8'd136;
	sample_rom[184][52] = 8'd130;
	sample_rom[184][53] = 8'd129;
	sample_rom[184][54] = 8'd129;
	sample_rom[184][55] = 8'd127;
	sample_rom[184][56] = 8'd129;
	sample_rom[184][57] = 8'd130;
	sample_rom[184][58] = 8'd132;
	sample_rom[184][59] = 8'd135;
	sample_rom[184][60] = 8'd136;
	sample_rom[184][61] = 8'd134;
	sample_rom[184][62] = 8'd131;
	sample_rom[184][63] = 8'd131;
	sample_rom[185][0] = 8'd131;
	sample_rom[185][1] = 8'd175;
	sample_rom[185][2] = 8'd211;
	sample_rom[185][3] = 8'd236;
	sample_rom[185][4] = 8'd250;
	sample_rom[185][5] = 8'd2;
	sample_rom[185][6] = 8'd246;
	sample_rom[185][7] = 8'd230;
	sample_rom[185][8] = 8'd211;
	sample_rom[185][9] = 8'd196;
	sample_rom[185][10] = 8'd183;
	sample_rom[185][11] = 8'd173;
	sample_rom[185][12] = 8'd172;
	sample_rom[185][13] = 8'd173;
	sample_rom[185][14] = 8'd178;
	sample_rom[185][15] = 8'd182;
	sample_rom[185][16] = 8'd185;
	sample_rom[185][17] = 8'd188;
	sample_rom[185][18] = 8'd186;
	sample_rom[185][19] = 8'd181;
	sample_rom[185][20] = 8'd177;
	sample_rom[185][21] = 8'd171;
	sample_rom[185][22] = 8'd166;
	sample_rom[185][23] = 8'd164;
	sample_rom[185][24] = 8'd165;
	sample_rom[185][25] = 8'd165;
	sample_rom[185][26] = 8'd165;
	sample_rom[185][27] = 8'd166;
	sample_rom[185][28] = 8'd165;
	sample_rom[185][29] = 8'd161;
	sample_rom[185][30] = 8'd159;
	sample_rom[185][31] = 8'd154;
	sample_rom[185][32] = 8'd151;
	sample_rom[185][33] = 8'd147;
	sample_rom[185][34] = 8'd149;
	sample_rom[185][35] = 8'd151;
	sample_rom[185][36] = 8'd150;
	sample_rom[185][37] = 8'd152;
	sample_rom[185][38] = 8'd153;
	sample_rom[185][39] = 8'd152;
	sample_rom[185][40] = 8'd153;
	sample_rom[185][41] = 8'd151;
	sample_rom[185][42] = 8'd147;
	sample_rom[185][43] = 8'd143;
	sample_rom[185][44] = 8'd140;
	sample_rom[185][45] = 8'd139;
	sample_rom[185][46] = 8'd138;
	sample_rom[185][47] = 8'd138;
	sample_rom[185][48] = 8'd140;
	sample_rom[185][49] = 8'd139;
	sample_rom[185][50] = 8'd139;
	sample_rom[185][51] = 8'd137;
	sample_rom[185][52] = 8'd135;
	sample_rom[185][53] = 8'd133;
	sample_rom[185][54] = 8'd130;
	sample_rom[185][55] = 8'd128;
	sample_rom[185][56] = 8'd126;
	sample_rom[185][57] = 8'd128;
	sample_rom[185][58] = 8'd129;
	sample_rom[185][59] = 8'd131;
	sample_rom[185][60] = 8'd131;
	sample_rom[185][61] = 8'd131;
	sample_rom[185][62] = 8'd130;
	sample_rom[185][63] = 8'd130;
	sample_rom[186][0] = 8'd130;
	sample_rom[186][1] = 8'd178;
	sample_rom[186][2] = 8'd217;
	sample_rom[186][3] = 8'd241;
	sample_rom[186][4] = 8'd252;
	sample_rom[186][5] = 8'd252;
	sample_rom[186][6] = 8'd238;
	sample_rom[186][7] = 8'd220;
	sample_rom[186][8] = 8'd199;
	sample_rom[186][9] = 8'd185;
	sample_rom[186][10] = 8'd174;
	sample_rom[186][11] = 8'd170;
	sample_rom[186][12] = 8'd173;
	sample_rom[186][13] = 8'd175;
	sample_rom[186][14] = 8'd180;
	sample_rom[186][15] = 8'd182;
	sample_rom[186][16] = 8'd182;
	sample_rom[186][17] = 8'd181;
	sample_rom[186][18] = 8'd176;
	sample_rom[186][19] = 8'd173;
	sample_rom[186][20] = 8'd170;
	sample_rom[186][21] = 8'd168;
	sample_rom[186][22] = 8'd171;
	sample_rom[186][23] = 8'd171;
	sample_rom[186][24] = 8'd173;
	sample_rom[186][25] = 8'd173;
	sample_rom[186][26] = 8'd170;
	sample_rom[186][27] = 8'd166;
	sample_rom[186][28] = 8'd162;
	sample_rom[186][29] = 8'd156;
	sample_rom[186][30] = 8'd155;
	sample_rom[186][31] = 8'd152;
	sample_rom[186][32] = 8'd153;
	sample_rom[186][33] = 8'd153;
	sample_rom[186][34] = 8'd158;
	sample_rom[186][35] = 8'd159;
	sample_rom[186][36] = 8'd156;
	sample_rom[186][37] = 8'd154;
	sample_rom[186][38] = 8'd150;
	sample_rom[186][39] = 8'd146;
	sample_rom[186][40] = 8'd145;
	sample_rom[186][41] = 8'd144;
	sample_rom[186][42] = 8'd143;
	sample_rom[186][43] = 8'd146;
	sample_rom[186][44] = 8'd145;
	sample_rom[186][45] = 8'd147;
	sample_rom[186][46] = 8'd145;
	sample_rom[186][47] = 8'd143;
	sample_rom[186][48] = 8'd140;
	sample_rom[186][49] = 8'd135;
	sample_rom[186][50] = 8'd131;
	sample_rom[186][51] = 8'd132;
	sample_rom[186][52] = 8'd131;
	sample_rom[186][53] = 8'd132;
	sample_rom[186][54] = 8'd135;
	sample_rom[186][55] = 8'd136;
	sample_rom[186][56] = 8'd135;
	sample_rom[186][57] = 8'd135;
	sample_rom[186][58] = 8'd134;
	sample_rom[186][59] = 8'd131;
	sample_rom[186][60] = 8'd126;
	sample_rom[186][61] = 8'd125;
	sample_rom[186][62] = 8'd124;
	sample_rom[186][63] = 8'd125;
	sample_rom[187][0] = 8'd130;
	sample_rom[187][1] = 8'd181;
	sample_rom[187][2] = 8'd223;
	sample_rom[187][3] = 8'd249;
	sample_rom[187][4] = 8'd3;
	sample_rom[187][5] = 8'd250;
	sample_rom[187][6] = 8'd234;
	sample_rom[187][7] = 8'd215;
	sample_rom[187][8] = 8'd195;
	sample_rom[187][9] = 8'd182;
	sample_rom[187][10] = 8'd176;
	sample_rom[187][11] = 8'd178;
	sample_rom[187][12] = 8'd184;
	sample_rom[187][13] = 8'd185;
	sample_rom[187][14] = 8'd189;
	sample_rom[187][15] = 8'd187;
	sample_rom[187][16] = 8'd185;
	sample_rom[187][17] = 8'd179;
	sample_rom[187][18] = 8'd174;
	sample_rom[187][19] = 8'd172;
	sample_rom[187][20] = 8'd168;
	sample_rom[187][21] = 8'd172;
	sample_rom[187][22] = 8'd172;
	sample_rom[187][23] = 8'd173;
	sample_rom[187][24] = 8'd171;
	sample_rom[187][25] = 8'd168;
	sample_rom[187][26] = 8'd162;
	sample_rom[187][27] = 8'd158;
	sample_rom[187][28] = 8'd155;
	sample_rom[187][29] = 8'd156;
	sample_rom[187][30] = 8'd158;
	sample_rom[187][31] = 8'd158;
	sample_rom[187][32] = 8'd160;
	sample_rom[187][33] = 8'd160;
	sample_rom[187][34] = 8'd160;
	sample_rom[187][35] = 8'd158;
	sample_rom[187][36] = 8'd152;
	sample_rom[187][37] = 8'd148;
	sample_rom[187][38] = 8'd146;
	sample_rom[187][39] = 8'd143;
	sample_rom[187][40] = 8'd145;
	sample_rom[187][41] = 8'd147;
	sample_rom[187][42] = 8'd147;
	sample_rom[187][43] = 8'd146;
	sample_rom[187][44] = 8'd144;
	sample_rom[187][45] = 8'd141;
	sample_rom[187][46] = 8'd138;
	sample_rom[187][47] = 8'd135;
	sample_rom[187][48] = 8'd133;
	sample_rom[187][49] = 8'd135;
	sample_rom[187][50] = 8'd136;
	sample_rom[187][51] = 8'd135;
	sample_rom[187][52] = 8'd137;
	sample_rom[187][53] = 8'd137;
	sample_rom[187][54] = 8'd134;
	sample_rom[187][55] = 8'd131;
	sample_rom[187][56] = 8'd131;
	sample_rom[187][57] = 8'd128;
	sample_rom[187][58] = 8'd129;
	sample_rom[187][59] = 8'd129;
	sample_rom[187][60] = 8'd129;
	sample_rom[187][61] = 8'd130;
	sample_rom[187][62] = 8'd130;
	sample_rom[187][63] = 8'd131;
	sample_rom[188][0] = 8'd130;
	sample_rom[188][1] = 8'd188;
	sample_rom[188][2] = 8'd228;
	sample_rom[188][3] = 8'd252;
	sample_rom[188][4] = 8'd253;
	sample_rom[188][5] = 8'd241;
	sample_rom[188][6] = 8'd220;
	sample_rom[188][7] = 8'd200;
	sample_rom[188][8] = 8'd185;
	sample_rom[188][9] = 8'd178;
	sample_rom[188][10] = 8'd179;
	sample_rom[188][11] = 8'd185;
	sample_rom[188][12] = 8'd188;
	sample_rom[188][13] = 8'd186;
	sample_rom[188][14] = 8'd185;
	sample_rom[188][15] = 8'd179;
	sample_rom[188][16] = 8'd175;
	sample_rom[188][17] = 8'd175;
	sample_rom[188][18] = 8'd175;
	sample_rom[188][19] = 8'd180;
	sample_rom[188][20] = 8'd178;
	sample_rom[188][21] = 8'd178;
	sample_rom[188][22] = 8'd175;
	sample_rom[188][23] = 8'd169;
	sample_rom[188][24] = 8'd165;
	sample_rom[188][25] = 8'd161;
	sample_rom[188][26] = 8'd161;
	sample_rom[188][27] = 8'd160;
	sample_rom[188][28] = 8'd161;
	sample_rom[188][29] = 8'd162;
	sample_rom[188][30] = 8'd163;
	sample_rom[188][31] = 8'd158;
	sample_rom[188][32] = 8'd154;
	sample_rom[188][33] = 8'd153;
	sample_rom[188][34] = 8'd151;
	sample_rom[188][35] = 8'd153;
	sample_rom[188][36] = 8'd150;
	sample_rom[188][37] = 8'd151;
	sample_rom[188][38] = 8'd150;
	sample_rom[188][39] = 8'd146;
	sample_rom[188][40] = 8'd145;
	sample_rom[188][41] = 8'd143;
	sample_rom[188][42] = 8'd145;
	sample_rom[188][43] = 8'd145;
	sample_rom[188][44] = 8'd146;
	sample_rom[188][45] = 8'd147;
	sample_rom[188][46] = 8'd146;
	sample_rom[188][47] = 8'd145;
	sample_rom[188][48] = 8'd140;
	sample_rom[188][49] = 8'd139;
	sample_rom[188][50] = 8'd136;
	sample_rom[188][51] = 8'd133;
	sample_rom[188][52] = 8'd136;
	sample_rom[188][53] = 8'd137;
	sample_rom[188][54] = 8'd135;
	sample_rom[188][55] = 8'd134;
	sample_rom[188][56] = 8'd134;
	sample_rom[188][57] = 8'd132;
	sample_rom[188][58] = 8'd133;
	sample_rom[188][59] = 8'd131;
	sample_rom[188][60] = 8'd128;
	sample_rom[188][61] = 8'd130;
	sample_rom[188][62] = 8'd129;
	sample_rom[188][63] = 8'd130;
	sample_rom[189][0] = 8'd130;
	sample_rom[189][1] = 8'd194;
	sample_rom[189][2] = 8'd239;
	sample_rom[189][3] = 8'd4;
	sample_rom[189][4] = 8'd246;
	sample_rom[189][5] = 8'd225;
	sample_rom[189][6] = 8'd201;
	sample_rom[189][7] = 8'd187;
	sample_rom[189][8] = 8'd181;
	sample_rom[189][9] = 8'd186;
	sample_rom[189][10] = 8'd189;
	sample_rom[189][11] = 8'd190;
	sample_rom[189][12] = 8'd183;
	sample_rom[189][13] = 8'd174;
	sample_rom[189][14] = 8'd171;
	sample_rom[189][15] = 8'd170;
	sample_rom[189][16] = 8'd173;
	sample_rom[189][17] = 8'd178;
	sample_rom[189][18] = 8'd180;
	sample_rom[189][19] = 8'd177;
	sample_rom[189][20] = 8'd169;
	sample_rom[189][21] = 8'd162;
	sample_rom[189][22] = 8'd160;
	sample_rom[189][23] = 8'd163;
	sample_rom[189][24] = 8'd167;
	sample_rom[189][25] = 8'd168;
	sample_rom[189][26] = 8'd170;
	sample_rom[189][27] = 8'd164;
	sample_rom[189][28] = 8'd157;
	sample_rom[189][29] = 8'd156;
	sample_rom[189][30] = 8'd154;
	sample_rom[189][31] = 8'd157;
	sample_rom[189][32] = 8'd157;
	sample_rom[189][33] = 8'd160;
	sample_rom[189][34] = 8'd156;
	sample_rom[189][35] = 8'd154;
	sample_rom[189][36] = 8'd149;
	sample_rom[189][37] = 8'd147;
	sample_rom[189][38] = 8'd149;
	sample_rom[189][39] = 8'd149;
	sample_rom[189][40] = 8'd150;
	sample_rom[189][41] = 8'd149;
	sample_rom[189][42] = 8'd146;
	sample_rom[189][43] = 8'd142;
	sample_rom[189][44] = 8'd141;
	sample_rom[189][45] = 8'd141;
	sample_rom[189][46] = 8'd143;
	sample_rom[189][47] = 8'd145;
	sample_rom[189][48] = 8'd144;
	sample_rom[189][49] = 8'd140;
	sample_rom[189][50] = 8'd137;
	sample_rom[189][51] = 8'd132;
	sample_rom[189][52] = 8'd136;
	sample_rom[189][53] = 8'd137;
	sample_rom[189][54] = 8'd137;
	sample_rom[189][55] = 8'd136;
	sample_rom[189][56] = 8'd137;
	sample_rom[189][57] = 8'd130;
	sample_rom[189][58] = 8'd127;
	sample_rom[189][59] = 8'd125;
	sample_rom[189][60] = 8'd123;
	sample_rom[189][61] = 8'd129;
	sample_rom[189][62] = 8'd129;
	sample_rom[189][63] = 8'd129;
	sample_rom[190][0] = 8'd130;
	sample_rom[190][1] = 8'd194;
	sample_rom[190][2] = 8'd235;
	sample_rom[190][3] = 8'd251;
	sample_rom[190][4] = 8'd242;
	sample_rom[190][5] = 8'd223;
	sample_rom[190][6] = 8'd200;
	sample_rom[190][7] = 8'd187;
	sample_rom[190][8] = 8'd183;
	sample_rom[190][9] = 8'd184;
	sample_rom[190][10] = 8'd183;
	sample_rom[190][11] = 8'd186;
	sample_rom[190][12] = 8'd179;
	sample_rom[190][13] = 8'd175;
	sample_rom[190][14] = 8'd177;
	sample_rom[190][15] = 8'd179;
	sample_rom[190][16] = 8'd179;
	sample_rom[190][17] = 8'd180;
	sample_rom[190][18] = 8'd177;
	sample_rom[190][19] = 8'd172;
	sample_rom[190][20] = 8'd170;
	sample_rom[190][21] = 8'd168;
	sample_rom[190][22] = 8'd168;
	sample_rom[190][23] = 8'd167;
	sample_rom[190][24] = 8'd167;
	sample_rom[190][25] = 8'd162;
	sample_rom[190][26] = 8'd161;
	sample_rom[190][27] = 8'd158;
	sample_rom[190][28] = 8'd156;
	sample_rom[190][29] = 8'd158;
	sample_rom[190][30] = 8'd157;
	sample_rom[190][31] = 8'd155;
	sample_rom[190][32] = 8'd154;
	sample_rom[190][33] = 8'd155;
	sample_rom[190][34] = 8'd153;
	sample_rom[190][35] = 8'd153;
	sample_rom[190][36] = 8'd152;
	sample_rom[190][37] = 8'd150;
	sample_rom[190][38] = 8'd152;
	sample_rom[190][39] = 8'd150;
	sample_rom[190][40] = 8'd149;
	sample_rom[190][41] = 8'd149;
	sample_rom[190][42] = 8'd148;
	sample_rom[190][43] = 8'd146;
	sample_rom[190][44] = 8'd145;
	sample_rom[190][45] = 8'd141;
	sample_rom[190][46] = 8'd141;
	sample_rom[190][47] = 8'd142;
	sample_rom[190][48] = 8'd143;
	sample_rom[190][49] = 8'd141;
	sample_rom[190][50] = 8'd136;
	sample_rom[190][51] = 8'd134;
	sample_rom[190][52] = 8'd135;
	sample_rom[190][53] = 8'd134;
	sample_rom[190][54] = 8'd133;
	sample_rom[190][55] = 8'd134;
	sample_rom[190][56] = 8'd138;
	sample_rom[190][57] = 8'd132;
	sample_rom[190][58] = 8'd129;
	sample_rom[190][59] = 8'd128;
	sample_rom[190][60] = 8'd123;
	sample_rom[190][61] = 8'd126;
	sample_rom[190][62] = 8'd127;
	sample_rom[190][63] = 8'd129;
	sample_rom[191][0] = 8'd130;
	sample_rom[191][1] = 8'd211;
	sample_rom[191][2] = 8'd4;
	sample_rom[191][3] = 8'd252;
	sample_rom[191][4] = 8'd223;
	sample_rom[191][5] = 8'd194;
	sample_rom[191][6] = 8'd183;
	sample_rom[191][7] = 8'd192;
	sample_rom[191][8] = 8'd197;
	sample_rom[191][9] = 8'd194;
	sample_rom[191][10] = 8'd179;
	sample_rom[191][11] = 8'd172;
	sample_rom[191][12] = 8'd168;
	sample_rom[191][13] = 8'd176;
	sample_rom[191][14] = 8'd181;
	sample_rom[191][15] = 8'd180;
	sample_rom[191][16] = 8'd174;
	sample_rom[191][17] = 8'd172;
	sample_rom[191][18] = 8'd175;
	sample_rom[191][19] = 8'd176;
	sample_rom[191][20] = 8'd175;
	sample_rom[191][21] = 8'd169;
	sample_rom[191][22] = 8'd164;
	sample_rom[191][23] = 8'd168;
	sample_rom[191][24] = 8'd172;
	sample_rom[191][25] = 8'd169;
	sample_rom[191][26] = 8'd170;
	sample_rom[191][27] = 8'd161;
	sample_rom[191][28] = 8'd157;
	sample_rom[191][29] = 8'd159;
	sample_rom[191][30] = 8'd159;
	sample_rom[191][31] = 8'd160;
	sample_rom[191][32] = 8'd156;
	sample_rom[191][33] = 8'd152;
	sample_rom[191][34] = 8'd149;
	sample_rom[191][35] = 8'd153;
	sample_rom[191][36] = 8'd157;
	sample_rom[191][37] = 8'd155;
	sample_rom[191][38] = 8'd154;
	sample_rom[191][39] = 8'd140;
	sample_rom[191][40] = 8'd141;
	sample_rom[191][41] = 8'd146;
	sample_rom[191][42] = 8'd150;
	sample_rom[191][43] = 8'd150;
	sample_rom[191][44] = 8'd146;
	sample_rom[191][45] = 8'd139;
	sample_rom[191][46] = 8'd141;
	sample_rom[191][47] = 8'd142;
	sample_rom[191][48] = 8'd145;
	sample_rom[191][49] = 8'd141;
	sample_rom[191][50] = 8'd137;
	sample_rom[191][51] = 8'd127;
	sample_rom[191][52] = 8'd130;
	sample_rom[191][53] = 8'd134;
	sample_rom[191][54] = 8'd136;
	sample_rom[191][55] = 8'd132;
	sample_rom[191][56] = 8'd133;
	sample_rom[191][57] = 8'd129;
	sample_rom[191][58] = 8'd131;
	sample_rom[191][59] = 8'd134;
	sample_rom[191][60] = 8'd132;
	sample_rom[191][61] = 8'd130;
	sample_rom[191][62] = 8'd125;
	sample_rom[191][63] = 8'd128;
	sample_rom[192][0] = 8'd130;
	sample_rom[192][1] = 8'd200;
	sample_rom[192][2] = 8'd237;
	sample_rom[192][3] = 8'd242;
	sample_rom[192][4] = 8'd224;
	sample_rom[192][5] = 8'd208;
	sample_rom[192][6] = 8'd192;
	sample_rom[192][7] = 8'd189;
	sample_rom[192][8] = 8'd185;
	sample_rom[192][9] = 8'd179;
	sample_rom[192][10] = 8'd175;
	sample_rom[192][11] = 8'd181;
	sample_rom[192][12] = 8'd182;
	sample_rom[192][13] = 8'd180;
	sample_rom[192][14] = 8'd177;
	sample_rom[192][15] = 8'd172;
	sample_rom[192][16] = 8'd172;
	sample_rom[192][17] = 8'd175;
	sample_rom[192][18] = 8'd176;
	sample_rom[192][19] = 8'd173;
	sample_rom[192][20] = 8'd169;
	sample_rom[192][21] = 8'd166;
	sample_rom[192][22] = 8'd165;
	sample_rom[192][23] = 8'd166;
	sample_rom[192][24] = 8'd168;
	sample_rom[192][25] = 8'd163;
	sample_rom[192][26] = 8'd162;
	sample_rom[192][27] = 8'd160;
	sample_rom[192][28] = 8'd158;
	sample_rom[192][29] = 8'd160;
	sample_rom[192][30] = 8'd158;
	sample_rom[192][31] = 8'd157;
	sample_rom[192][32] = 8'd157;
	sample_rom[192][33] = 8'd159;
	sample_rom[192][34] = 8'd155;
	sample_rom[192][35] = 8'd151;
	sample_rom[192][36] = 8'd149;
	sample_rom[192][37] = 8'd144;
	sample_rom[192][38] = 8'd149;
	sample_rom[192][39] = 8'd145;
	sample_rom[192][40] = 8'd145;
	sample_rom[192][41] = 8'd142;
	sample_rom[192][42] = 8'd141;
	sample_rom[192][43] = 8'd142;
	sample_rom[192][44] = 8'd144;
	sample_rom[192][45] = 8'd140;
	sample_rom[192][46] = 8'd142;
	sample_rom[192][47] = 8'd143;
	sample_rom[192][48] = 8'd143;
	sample_rom[192][49] = 8'd140;
	sample_rom[192][50] = 8'd137;
	sample_rom[192][51] = 8'd133;
	sample_rom[192][52] = 8'd131;
	sample_rom[192][53] = 8'd130;
	sample_rom[192][54] = 8'd132;
	sample_rom[192][55] = 8'd132;
	sample_rom[192][56] = 8'd134;
	sample_rom[192][57] = 8'd130;
	sample_rom[192][58] = 8'd131;
	sample_rom[192][59] = 8'd131;
	sample_rom[192][60] = 8'd127;
	sample_rom[192][61] = 8'd128;
	sample_rom[192][62] = 8'd127;
	sample_rom[192][63] = 8'd129;
	sample_rom[193][0] = 8'd130;
	sample_rom[193][1] = 8'd217;
	sample_rom[193][2] = 8'd4;
	sample_rom[193][3] = 8'd245;
	sample_rom[193][4] = 8'd208;
	sample_rom[193][5] = 8'd178;
	sample_rom[193][6] = 8'd176;
	sample_rom[193][7] = 8'd193;
	sample_rom[193][8] = 8'd203;
	sample_rom[193][9] = 8'd197;
	sample_rom[193][10] = 8'd184;
	sample_rom[193][11] = 8'd172;
	sample_rom[193][12] = 8'd173;
	sample_rom[193][13] = 8'd179;
	sample_rom[193][14] = 8'd177;
	sample_rom[193][15] = 8'd175;
	sample_rom[193][16] = 8'd171;
	sample_rom[193][17] = 8'd173;
	sample_rom[193][18] = 8'd179;
	sample_rom[193][19] = 8'd181;
	sample_rom[193][20] = 8'd177;
	sample_rom[193][21] = 8'd168;
	sample_rom[193][22] = 8'd159;
	sample_rom[193][23] = 8'd161;
	sample_rom[193][24] = 8'd163;
	sample_rom[193][25] = 8'd165;
	sample_rom[193][26] = 8'd164;
	sample_rom[193][27] = 8'd163;
	sample_rom[193][28] = 8'd160;
	sample_rom[193][29] = 8'd157;
	sample_rom[193][30] = 8'd157;
	sample_rom[193][31] = 8'd156;
	sample_rom[193][32] = 8'd155;
	sample_rom[193][33] = 8'd156;
	sample_rom[193][34] = 8'd150;
	sample_rom[193][35] = 8'd152;
	sample_rom[193][36] = 8'd153;
	sample_rom[193][37] = 8'd149;
	sample_rom[193][38] = 8'd152;
	sample_rom[193][39] = 8'd143;
	sample_rom[193][40] = 8'd143;
	sample_rom[193][41] = 8'd143;
	sample_rom[193][42] = 8'd147;
	sample_rom[193][43] = 8'd146;
	sample_rom[193][44] = 8'd143;
	sample_rom[193][45] = 8'd137;
	sample_rom[193][46] = 8'd135;
	sample_rom[193][47] = 8'd134;
	sample_rom[193][48] = 8'd135;
	sample_rom[193][49] = 8'd136;
	sample_rom[193][50] = 8'd138;
	sample_rom[193][51] = 8'd131;
	sample_rom[193][52] = 8'd134;
	sample_rom[193][53] = 8'd137;
	sample_rom[193][54] = 8'd139;
	sample_rom[193][55] = 8'd134;
	sample_rom[193][56] = 8'd131;
	sample_rom[193][57] = 8'd129;
	sample_rom[193][58] = 8'd130;
	sample_rom[193][59] = 8'd132;
	sample_rom[193][60] = 8'd131;
	sample_rom[193][61] = 8'd128;
	sample_rom[193][62] = 8'd126;
	sample_rom[193][63] = 8'd127;
	sample_rom[194][0] = 8'd130;
	sample_rom[194][1] = 8'd195;
	sample_rom[194][2] = 8'd227;
	sample_rom[194][3] = 8'd231;
	sample_rom[194][4] = 8'd213;
	sample_rom[194][5] = 8'd197;
	sample_rom[194][6] = 8'd184;
	sample_rom[194][7] = 8'd184;
	sample_rom[194][8] = 8'd185;
	sample_rom[194][9] = 8'd178;
	sample_rom[194][10] = 8'd177;
	sample_rom[194][11] = 8'd178;
	sample_rom[194][12] = 8'd181;
	sample_rom[194][13] = 8'd179;
	sample_rom[194][14] = 8'd176;
	sample_rom[194][15] = 8'd171;
	sample_rom[194][16] = 8'd171;
	sample_rom[194][17] = 8'd174;
	sample_rom[194][18] = 8'd177;
	sample_rom[194][19] = 8'd174;
	sample_rom[194][20] = 8'd172;
	sample_rom[194][21] = 8'd166;
	sample_rom[194][22] = 8'd165;
	sample_rom[194][23] = 8'd168;
	sample_rom[194][24] = 8'd167;
	sample_rom[194][25] = 8'd164;
	sample_rom[194][26] = 8'd160;
	sample_rom[194][27] = 8'd161;
	sample_rom[194][28] = 8'd159;
	sample_rom[194][29] = 8'd159;
	sample_rom[194][30] = 8'd160;
	sample_rom[194][31] = 8'd156;
	sample_rom[194][32] = 8'd155;
	sample_rom[194][33] = 8'd155;
	sample_rom[194][34] = 8'd151;
	sample_rom[194][35] = 8'd147;
	sample_rom[194][36] = 8'd145;
	sample_rom[194][37] = 8'd142;
	sample_rom[194][38] = 8'd150;
	sample_rom[194][39] = 8'd148;
	sample_rom[194][40] = 8'd150;
	sample_rom[194][41] = 8'd146;
	sample_rom[194][42] = 8'd147;
	sample_rom[194][43] = 8'd144;
	sample_rom[194][44] = 8'd145;
	sample_rom[194][45] = 8'd142;
	sample_rom[194][46] = 8'd142;
	sample_rom[194][47] = 8'd142;
	sample_rom[194][48] = 8'd140;
	sample_rom[194][49] = 8'd138;
	sample_rom[194][50] = 8'd138;
	sample_rom[194][51] = 8'd134;
	sample_rom[194][52] = 8'd134;
	sample_rom[194][53] = 8'd133;
	sample_rom[194][54] = 8'd134;
	sample_rom[194][55] = 8'd138;
	sample_rom[194][56] = 8'd135;
	sample_rom[194][57] = 8'd134;
	sample_rom[194][58] = 8'd135;
	sample_rom[194][59] = 8'd134;
	sample_rom[194][60] = 8'd131;
	sample_rom[194][61] = 8'd129;
	sample_rom[194][62] = 8'd129;
	sample_rom[194][63] = 8'd128;
	sample_rom[195][0] = 8'd130;
	sample_rom[195][1] = 8'd208;
	sample_rom[195][2] = 8'd252;
	sample_rom[195][3] = 8'd4;
	sample_rom[195][4] = 8'd233;
	sample_rom[195][5] = 8'd214;
	sample_rom[195][6] = 8'd199;
	sample_rom[195][7] = 8'd198;
	sample_rom[195][8] = 8'd194;
	sample_rom[195][9] = 8'd192;
	sample_rom[195][10] = 8'd190;
	sample_rom[195][11] = 8'd192;
	sample_rom[195][12] = 8'd191;
	sample_rom[195][13] = 8'd181;
	sample_rom[195][14] = 8'd177;
	sample_rom[195][15] = 8'd169;
	sample_rom[195][16] = 8'd170;
	sample_rom[195][17] = 8'd175;
	sample_rom[195][18] = 8'd180;
	sample_rom[195][19] = 8'd176;
	sample_rom[195][20] = 8'd169;
	sample_rom[195][21] = 8'd163;
	sample_rom[195][22] = 8'd163;
	sample_rom[195][23] = 8'd166;
	sample_rom[195][24] = 8'd165;
	sample_rom[195][25] = 8'd163;
	sample_rom[195][26] = 8'd163;
	sample_rom[195][27] = 8'd160;
	sample_rom[195][28] = 8'd154;
	sample_rom[195][29] = 8'd157;
	sample_rom[195][30] = 8'd154;
	sample_rom[195][31] = 8'd151;
	sample_rom[195][32] = 8'd150;
	sample_rom[195][33] = 8'd153;
	sample_rom[195][34] = 8'd148;
	sample_rom[195][35] = 8'd145;
	sample_rom[195][36] = 8'd142;
	sample_rom[195][37] = 8'd138;
	sample_rom[195][38] = 8'd143;
	sample_rom[195][39] = 8'd141;
	sample_rom[195][40] = 8'd143;
	sample_rom[195][41] = 8'd141;
	sample_rom[195][42] = 8'd138;
	sample_rom[195][43] = 8'd136;
	sample_rom[195][44] = 8'd137;
	sample_rom[195][45] = 8'd137;
	sample_rom[195][46] = 8'd141;
	sample_rom[195][47] = 8'd142;
	sample_rom[195][48] = 8'd141;
	sample_rom[195][49] = 8'd139;
	sample_rom[195][50] = 8'd133;
	sample_rom[195][51] = 8'd127;
	sample_rom[195][52] = 8'd128;
	sample_rom[195][53] = 8'd128;
	sample_rom[195][54] = 8'd131;
	sample_rom[195][55] = 8'd131;
	sample_rom[195][56] = 8'd135;
	sample_rom[195][57] = 8'd129;
	sample_rom[195][58] = 8'd130;
	sample_rom[195][59] = 8'd129;
	sample_rom[195][60] = 8'd126;
	sample_rom[195][61] = 8'd131;
	sample_rom[195][62] = 8'd129;
	sample_rom[195][63] = 8'd130;
	sample_rom[196][0] = 8'd130;
	sample_rom[196][1] = 8'd189;
	sample_rom[196][2] = 8'd220;
	sample_rom[196][3] = 8'd223;
	sample_rom[196][4] = 8'd206;
	sample_rom[196][5] = 8'd193;
	sample_rom[196][6] = 8'd184;
	sample_rom[196][7] = 8'd185;
	sample_rom[196][8] = 8'd186;
	sample_rom[196][9] = 8'd177;
	sample_rom[196][10] = 8'd174;
	sample_rom[196][11] = 8'd174;
	sample_rom[196][12] = 8'd177;
	sample_rom[196][13] = 8'd173;
	sample_rom[196][14] = 8'd173;
	sample_rom[196][15] = 8'd168;
	sample_rom[196][16] = 8'd169;
	sample_rom[196][17] = 8'd172;
	sample_rom[196][18] = 8'd174;
	sample_rom[196][19] = 8'd167;
	sample_rom[196][20] = 8'd165;
	sample_rom[196][21] = 8'd160;
	sample_rom[196][22] = 8'd160;
	sample_rom[196][23] = 8'd165;
	sample_rom[196][24] = 8'd163;
	sample_rom[196][25] = 8'd163;
	sample_rom[196][26] = 8'd158;
	sample_rom[196][27] = 8'd160;
	sample_rom[196][28] = 8'd157;
	sample_rom[196][29] = 8'd155;
	sample_rom[196][30] = 8'd156;
	sample_rom[196][31] = 8'd152;
	sample_rom[196][32] = 8'd153;
	sample_rom[196][33] = 8'd155;
	sample_rom[196][34] = 8'd152;
	sample_rom[196][35] = 8'd151;
	sample_rom[196][36] = 8'd148;
	sample_rom[196][37] = 8'd140;
	sample_rom[196][38] = 8'd145;
	sample_rom[196][39] = 8'd142;
	sample_rom[196][40] = 8'd142;
	sample_rom[196][41] = 8'd138;
	sample_rom[196][42] = 8'd138;
	sample_rom[196][43] = 8'd137;
	sample_rom[196][44] = 8'd141;
	sample_rom[196][45] = 8'd140;
	sample_rom[196][46] = 8'd141;
	sample_rom[196][47] = 8'd140;
	sample_rom[196][48] = 8'd138;
	sample_rom[196][49] = 8'd138;
	sample_rom[196][50] = 8'd135;
	sample_rom[196][51] = 8'd133;
	sample_rom[196][52] = 8'd130;
	sample_rom[196][53] = 8'd130;
	sample_rom[196][54] = 8'd130;
	sample_rom[196][55] = 8'd133;
	sample_rom[196][56] = 8'd130;
	sample_rom[196][57] = 8'd129;
	sample_rom[196][58] = 8'd131;
	sample_rom[196][59] = 8'd130;
	sample_rom[196][60] = 8'd129;
	sample_rom[196][61] = 8'd128;
	sample_rom[196][62] = 8'd129;
	sample_rom[196][63] = 8'd128;
	sample_rom[197][0] = 8'd130;
	sample_rom[197][1] = 8'd204;
	sample_rom[197][2] = 8'd252;
	sample_rom[197][3] = 8'd13;
	sample_rom[197][4] = 8'd251;
	sample_rom[197][5] = 8'd233;
	sample_rom[197][6] = 8'd222;
	sample_rom[197][7] = 8'd215;
	sample_rom[197][8] = 8'd213;
	sample_rom[197][9] = 8'd211;
	sample_rom[197][10] = 8'd210;
	sample_rom[197][11] = 8'd208;
	sample_rom[197][12] = 8'd208;
	sample_rom[197][13] = 8'd203;
	sample_rom[197][14] = 8'd198;
	sample_rom[197][15] = 8'd196;
	sample_rom[197][16] = 8'd195;
	sample_rom[197][17] = 8'd196;
	sample_rom[197][18] = 8'd198;
	sample_rom[197][19] = 8'd191;
	sample_rom[197][20] = 8'd185;
	sample_rom[197][21] = 8'd182;
	sample_rom[197][22] = 8'd181;
	sample_rom[197][23] = 8'd185;
	sample_rom[197][24] = 8'd178;
	sample_rom[197][25] = 8'd178;
	sample_rom[197][26] = 8'd175;
	sample_rom[197][27] = 8'd174;
	sample_rom[197][28] = 8'd169;
	sample_rom[197][29] = 8'd169;
	sample_rom[197][30] = 8'd166;
	sample_rom[197][31] = 8'd164;
	sample_rom[197][32] = 8'd163;
	sample_rom[197][33] = 8'd161;
	sample_rom[197][34] = 8'd161;
	sample_rom[197][35] = 8'd158;
	sample_rom[197][36] = 8'd154;
	sample_rom[197][37] = 8'd155;
	sample_rom[197][38] = 8'd157;
	sample_rom[197][39] = 8'd155;
	sample_rom[197][40] = 8'd153;
	sample_rom[197][41] = 8'd147;
	sample_rom[197][42] = 8'd147;
	sample_rom[197][43] = 8'd145;
	sample_rom[197][44] = 8'd144;
	sample_rom[197][45] = 8'd141;
	sample_rom[197][46] = 8'd140;
	sample_rom[197][47] = 8'd138;
	sample_rom[197][48] = 8'd138;
	sample_rom[197][49] = 8'd136;
	sample_rom[197][50] = 8'd135;
	sample_rom[197][51] = 8'd129;
	sample_rom[197][52] = 8'd130;
	sample_rom[197][53] = 8'd133;
	sample_rom[197][54] = 8'd135;
	sample_rom[197][55] = 8'd133;
	sample_rom[197][56] = 8'd132;
	sample_rom[197][57] = 8'd132;
	sample_rom[197][58] = 8'd133;
	sample_rom[197][59] = 8'd131;
	sample_rom[197][60] = 8'd130;
	sample_rom[197][61] = 8'd131;
	sample_rom[197][62] = 8'd126;
	sample_rom[197][63] = 8'd127;
	sample_rom[198][0] = 8'd130;
	sample_rom[198][1] = 8'd184;
	sample_rom[198][2] = 8'd212;
	sample_rom[198][3] = 8'd214;
	sample_rom[198][4] = 8'd196;
	sample_rom[198][5] = 8'd187;
	sample_rom[198][6] = 8'd182;
	sample_rom[198][7] = 8'd183;
	sample_rom[198][8] = 8'd180;
	sample_rom[198][9] = 8'd175;
	sample_rom[198][10] = 8'd170;
	sample_rom[198][11] = 8'd170;
	sample_rom[198][12] = 8'd174;
	sample_rom[198][13] = 8'd171;
	sample_rom[198][14] = 8'd172;
	sample_rom[198][15] = 8'd165;
	sample_rom[198][16] = 8'd166;
	sample_rom[198][17] = 8'd168;
	sample_rom[198][18] = 8'd170;
	sample_rom[198][19] = 8'd162;
	sample_rom[198][20] = 8'd162;
	sample_rom[198][21] = 8'd158;
	sample_rom[198][22] = 8'd159;
	sample_rom[198][23] = 8'd164;
	sample_rom[198][24] = 8'd161;
	sample_rom[198][25] = 8'd158;
	sample_rom[198][26] = 8'd153;
	sample_rom[198][27] = 8'd152;
	sample_rom[198][28] = 8'd146;
	sample_rom[198][29] = 8'd149;
	sample_rom[198][30] = 8'd149;
	sample_rom[198][31] = 8'd148;
	sample_rom[198][32] = 8'd149;
	sample_rom[198][33] = 8'd152;
	sample_rom[198][34] = 8'd150;
	sample_rom[198][35] = 8'd145;
	sample_rom[198][36] = 8'd144;
	sample_rom[198][37] = 8'd138;
	sample_rom[198][38] = 8'd144;
	sample_rom[198][39] = 8'd143;
	sample_rom[198][40] = 8'd146;
	sample_rom[198][41] = 8'd142;
	sample_rom[198][42] = 8'd141;
	sample_rom[198][43] = 8'd138;
	sample_rom[198][44] = 8'd138;
	sample_rom[198][45] = 8'd137;
	sample_rom[198][46] = 8'd137;
	sample_rom[198][47] = 8'd136;
	sample_rom[198][48] = 8'd137;
	sample_rom[198][49] = 8'd136;
	sample_rom[198][50] = 8'd133;
	sample_rom[198][51] = 8'd132;
	sample_rom[198][52] = 8'd129;
	sample_rom[198][53] = 8'd130;
	sample_rom[198][54] = 8'd131;
	sample_rom[198][55] = 8'd135;
	sample_rom[198][56] = 8'd132;
	sample_rom[198][57] = 8'd130;
	sample_rom[198][58] = 8'd131;
	sample_rom[198][59] = 8'd130;
	sample_rom[198][60] = 8'd123;
	sample_rom[198][61] = 8'd125;
	sample_rom[198][62] = 8'd123;
	sample_rom[198][63] = 8'd124;
	sample_rom[199][0] = 8'd130;
	sample_rom[199][1] = 8'd198;
	sample_rom[199][2] = 8'd244;
	sample_rom[199][3] = 8'd6;
	sample_rom[199][4] = 8'd250;
	sample_rom[199][5] = 8'd233;
	sample_rom[199][6] = 8'd223;
	sample_rom[199][7] = 8'd215;
	sample_rom[199][8] = 8'd209;
	sample_rom[199][9] = 8'd200;
	sample_rom[199][10] = 8'd195;
	sample_rom[199][11] = 8'd192;
	sample_rom[199][12] = 8'd196;
	sample_rom[199][13] = 8'd195;
	sample_rom[199][14] = 8'd195;
	sample_rom[199][15] = 8'd192;
	sample_rom[199][16] = 8'd190;
	sample_rom[199][17] = 8'd191;
	sample_rom[199][18] = 8'd193;
	sample_rom[199][19] = 8'd187;
	sample_rom[199][20] = 8'd182;
	sample_rom[199][21] = 8'd177;
	sample_rom[199][22] = 8'd180;
	sample_rom[199][23] = 8'd176;
	sample_rom[199][24] = 8'd171;
	sample_rom[199][25] = 8'd166;
	sample_rom[199][26] = 8'd162;
	sample_rom[199][27] = 8'd162;
	sample_rom[199][28] = 8'd159;
	sample_rom[199][29] = 8'd161;
	sample_rom[199][30] = 8'd160;
	sample_rom[199][31] = 8'd158;
	sample_rom[199][32] = 8'd157;
	sample_rom[199][33] = 8'd157;
	sample_rom[199][34] = 8'd153;
	sample_rom[199][35] = 8'd151;
	sample_rom[199][36] = 8'd148;
	sample_rom[199][37] = 8'd148;
	sample_rom[199][38] = 8'd153;
	sample_rom[199][39] = 8'd153;
	sample_rom[199][40] = 8'd150;
	sample_rom[199][41] = 8'd145;
	sample_rom[199][42] = 8'd144;
	sample_rom[199][43] = 8'd147;
	sample_rom[199][44] = 8'd144;
	sample_rom[199][45] = 8'd143;
	sample_rom[199][46] = 8'd141;
	sample_rom[199][47] = 8'd137;
	sample_rom[199][48] = 8'd139;
	sample_rom[199][49] = 8'd137;
	sample_rom[199][50] = 8'd139;
	sample_rom[199][51] = 8'd134;
	sample_rom[199][52] = 8'd132;
	sample_rom[199][53] = 8'd131;
	sample_rom[199][54] = 8'd133;
	sample_rom[199][55] = 8'd128;
	sample_rom[199][56] = 8'd125;
	sample_rom[199][57] = 8'd127;
	sample_rom[199][58] = 8'd127;
	sample_rom[199][59] = 8'd130;
	sample_rom[199][60] = 8'd129;
	sample_rom[199][61] = 8'd132;
	sample_rom[199][62] = 8'd125;
	sample_rom[199][63] = 8'd129;
	sample_rom[200][0] = 8'd130;
	sample_rom[200][1] = 8'd177;
	sample_rom[200][2] = 8'd203;
	sample_rom[200][3] = 8'd205;
	sample_rom[200][4] = 8'd192;
	sample_rom[200][5] = 8'd185;
	sample_rom[200][6] = 8'd182;
	sample_rom[200][7] = 8'd184;
	sample_rom[200][8] = 8'd178;
	sample_rom[200][9] = 8'd170;
	sample_rom[200][10] = 8'd166;
	sample_rom[200][11] = 8'd166;
	sample_rom[200][12] = 8'd172;
	sample_rom[200][13] = 8'd171;
	sample_rom[200][14] = 8'd172;
	sample_rom[200][15] = 8'd164;
	sample_rom[200][16] = 8'd161;
	sample_rom[200][17] = 8'd162;
	sample_rom[200][18] = 8'd164;
	sample_rom[200][19] = 8'd160;
	sample_rom[200][20] = 8'd160;
	sample_rom[200][21] = 8'd159;
	sample_rom[200][22] = 8'd159;
	sample_rom[200][23] = 8'd162;
	sample_rom[200][24] = 8'd156;
	sample_rom[200][25] = 8'd153;
	sample_rom[200][26] = 8'd149;
	sample_rom[200][27] = 8'd150;
	sample_rom[200][28] = 8'd149;
	sample_rom[200][29] = 8'd154;
	sample_rom[200][30] = 8'd151;
	sample_rom[200][31] = 8'd146;
	sample_rom[200][32] = 8'd143;
	sample_rom[200][33] = 8'd141;
	sample_rom[200][34] = 8'd140;
	sample_rom[200][35] = 8'd136;
	sample_rom[200][36] = 8'd138;
	sample_rom[200][37] = 8'd133;
	sample_rom[200][38] = 8'd140;
	sample_rom[200][39] = 8'd138;
	sample_rom[200][40] = 8'd141;
	sample_rom[200][41] = 8'd137;
	sample_rom[200][42] = 8'd138;
	sample_rom[200][43] = 8'd136;
	sample_rom[200][44] = 8'd136;
	sample_rom[200][45] = 8'd135;
	sample_rom[200][46] = 8'd133;
	sample_rom[200][47] = 8'd133;
	sample_rom[200][48] = 8'd132;
	sample_rom[200][49] = 8'd132;
	sample_rom[200][50] = 8'd130;
	sample_rom[200][51] = 8'd130;
	sample_rom[200][52] = 8'd128;
	sample_rom[200][53] = 8'd130;
	sample_rom[200][54] = 8'd131;
	sample_rom[200][55] = 8'd133;
	sample_rom[200][56] = 8'd131;
	sample_rom[200][57] = 8'd129;
	sample_rom[200][58] = 8'd132;
	sample_rom[200][59] = 8'd131;
	sample_rom[200][60] = 8'd127;
	sample_rom[200][61] = 8'd130;
	sample_rom[200][62] = 8'd127;
	sample_rom[200][63] = 8'd126;
	sample_rom[201][0] = 8'd131;
	sample_rom[201][1] = 8'd205;
	sample_rom[201][2] = 8'd245;
	sample_rom[201][3] = 8'd9;
	sample_rom[201][4] = 8'd248;
	sample_rom[201][5] = 8'd230;
	sample_rom[201][6] = 8'd224;
	sample_rom[201][7] = 8'd221;
	sample_rom[201][8] = 8'd216;
	sample_rom[201][9] = 8'd204;
	sample_rom[201][10] = 8'd198;
	sample_rom[201][11] = 8'd194;
	sample_rom[201][12] = 8'd196;
	sample_rom[201][13] = 8'd194;
	sample_rom[201][14] = 8'd193;
	sample_rom[201][15] = 8'd192;
	sample_rom[201][16] = 8'd192;
	sample_rom[201][17] = 8'd191;
	sample_rom[201][18] = 8'd188;
	sample_rom[201][19] = 8'd183;
	sample_rom[201][20] = 8'd178;
	sample_rom[201][21] = 8'd178;
	sample_rom[201][22] = 8'd178;
	sample_rom[201][23] = 8'd178;
	sample_rom[201][24] = 8'd172;
	sample_rom[201][25] = 8'd169;
	sample_rom[201][26] = 8'd160;
	sample_rom[201][27] = 8'd162;
	sample_rom[201][28] = 8'd160;
	sample_rom[201][29] = 8'd160;
	sample_rom[201][30] = 8'd160;
	sample_rom[201][31] = 8'd156;
	sample_rom[201][32] = 8'd152;
	sample_rom[201][33] = 8'd151;
	sample_rom[201][34] = 8'd150;
	sample_rom[201][35] = 8'd145;
	sample_rom[201][36] = 8'd148;
	sample_rom[201][37] = 8'd143;
	sample_rom[201][38] = 8'd142;
	sample_rom[201][39] = 8'd142;
	sample_rom[201][40] = 8'd140;
	sample_rom[201][41] = 8'd140;
	sample_rom[201][42] = 8'd138;
	sample_rom[201][43] = 8'd141;
	sample_rom[201][44] = 8'd140;
	sample_rom[201][45] = 8'd140;
	sample_rom[201][46] = 8'd138;
	sample_rom[201][47] = 8'd138;
	sample_rom[201][48] = 8'd138;
	sample_rom[201][49] = 8'd139;
	sample_rom[201][50] = 8'd138;
	sample_rom[201][51] = 8'd133;
	sample_rom[201][52] = 8'd130;
	sample_rom[201][53] = 8'd130;
	sample_rom[201][54] = 8'd134;
	sample_rom[201][55] = 8'd133;
	sample_rom[201][56] = 8'd135;
	sample_rom[201][57] = 8'd130;
	sample_rom[201][58] = 8'd131;
	sample_rom[201][59] = 8'd126;
	sample_rom[201][60] = 8'd128;
	sample_rom[201][61] = 8'd126;
	sample_rom[201][62] = 8'd127;
	sample_rom[201][63] = 8'd126;
	sample_rom[202][0] = 8'd129;
	sample_rom[202][1] = 8'd176;
	sample_rom[202][2] = 8'd200;
	sample_rom[202][3] = 8'd202;
	sample_rom[202][4] = 8'd190;
	sample_rom[202][5] = 8'd182;
	sample_rom[202][6] = 8'd180;
	sample_rom[202][7] = 8'd183;
	sample_rom[202][8] = 8'd176;
	sample_rom[202][9] = 8'd168;
	sample_rom[202][10] = 8'd164;
	sample_rom[202][11] = 8'd163;
	sample_rom[202][12] = 8'd169;
	sample_rom[202][13] = 8'd167;
	sample_rom[202][14] = 8'd167;
	sample_rom[202][15] = 8'd159;
	sample_rom[202][16] = 8'd155;
	sample_rom[202][17] = 8'd156;
	sample_rom[202][18] = 8'd159;
	sample_rom[202][19] = 8'd155;
	sample_rom[202][20] = 8'd157;
	sample_rom[202][21] = 8'd155;
	sample_rom[202][22] = 8'd157;
	sample_rom[202][23] = 8'd159;
	sample_rom[202][24] = 8'd152;
	sample_rom[202][25] = 8'd148;
	sample_rom[202][26] = 8'd144;
	sample_rom[202][27] = 8'd146;
	sample_rom[202][28] = 8'd143;
	sample_rom[202][29] = 8'd147;
	sample_rom[202][30] = 8'd144;
	sample_rom[202][31] = 8'd140;
	sample_rom[202][32] = 8'd140;
	sample_rom[202][33] = 8'd139;
	sample_rom[202][34] = 8'd139;
	sample_rom[202][35] = 8'd135;
	sample_rom[202][36] = 8'd137;
	sample_rom[202][37] = 8'd131;
	sample_rom[202][38] = 8'd137;
	sample_rom[202][39] = 8'd135;
	sample_rom[202][40] = 8'd137;
	sample_rom[202][41] = 8'd133;
	sample_rom[202][42] = 8'd134;
	sample_rom[202][43] = 8'd134;
	sample_rom[202][44] = 8'd134;
	sample_rom[202][45] = 8'd135;
	sample_rom[202][46] = 8'd133;
	sample_rom[202][47] = 8'd134;
	sample_rom[202][48] = 8'd134;
	sample_rom[202][49] = 8'd134;
	sample_rom[202][50] = 8'd131;
	sample_rom[202][51] = 8'd130;
	sample_rom[202][52] = 8'd128;
	sample_rom[202][53] = 8'd127;
	sample_rom[202][54] = 8'd128;
	sample_rom[202][55] = 8'd131;
	sample_rom[202][56] = 8'd131;
	sample_rom[202][57] = 8'd128;
	sample_rom[202][58] = 8'd132;
	sample_rom[202][59] = 8'd131;
	sample_rom[202][60] = 8'd129;
	sample_rom[202][61] = 8'd132;
	sample_rom[202][62] = 8'd130;
	sample_rom[202][63] = 8'd128;
	sample_rom[203][0] = 8'd131;
	sample_rom[203][1] = 8'd213;
	sample_rom[203][2] = 8'd253;
	sample_rom[203][3] = 8'd10;
	sample_rom[203][4] = 8'd240;
	sample_rom[203][5] = 8'd218;
	sample_rom[203][6] = 8'd206;
	sample_rom[203][7] = 8'd202;
	sample_rom[203][8] = 8'd199;
	sample_rom[203][9] = 8'd189;
	sample_rom[203][10] = 8'd183;
	sample_rom[203][11] = 8'd181;
	sample_rom[203][12] = 8'd180;
	sample_rom[203][13] = 8'd180;
	sample_rom[203][14] = 8'd176;
	sample_rom[203][15] = 8'd172;
	sample_rom[203][16] = 8'd167;
	sample_rom[203][17] = 8'd168;
	sample_rom[203][18] = 8'd168;
	sample_rom[203][19] = 8'd167;
	sample_rom[203][20] = 8'd165;
	sample_rom[203][21] = 8'd163;
	sample_rom[203][22] = 8'd160;
	sample_rom[203][23] = 8'd160;
	sample_rom[203][24] = 8'd157;
	sample_rom[203][25] = 8'd154;
	sample_rom[203][26] = 8'd151;
	sample_rom[203][27] = 8'd155;
	sample_rom[203][28] = 8'd151;
	sample_rom[203][29] = 8'd151;
	sample_rom[203][30] = 8'd147;
	sample_rom[203][31] = 8'd144;
	sample_rom[203][32] = 8'd143;
	sample_rom[203][33] = 8'd145;
	sample_rom[203][34] = 8'd145;
	sample_rom[203][35] = 8'd143;
	sample_rom[203][36] = 8'd142;
	sample_rom[203][37] = 8'd140;
	sample_rom[203][38] = 8'd141;
	sample_rom[203][39] = 8'd143;
	sample_rom[203][40] = 8'd140;
	sample_rom[203][41] = 8'd138;
	sample_rom[203][42] = 8'd138;
	sample_rom[203][43] = 8'd139;
	sample_rom[203][44] = 8'd138;
	sample_rom[203][45] = 8'd138;
	sample_rom[203][46] = 8'd136;
	sample_rom[203][47] = 8'd136;
	sample_rom[203][48] = 8'd137;
	sample_rom[203][49] = 8'd139;
	sample_rom[203][50] = 8'd138;
	sample_rom[203][51] = 8'd136;
	sample_rom[203][52] = 8'd133;
	sample_rom[203][53] = 8'd128;
	sample_rom[203][54] = 8'd129;
	sample_rom[203][55] = 8'd128;
	sample_rom[203][56] = 8'd131;
	sample_rom[203][57] = 8'd129;
	sample_rom[203][58] = 8'd130;
	sample_rom[203][59] = 8'd129;
	sample_rom[203][60] = 8'd127;
	sample_rom[203][61] = 8'd127;
	sample_rom[203][62] = 8'd128;
	sample_rom[203][63] = 8'd126;
	sample_rom[204][0] = 8'd128;
	sample_rom[204][1] = 8'd170;
	sample_rom[204][2] = 8'd194;
	sample_rom[204][3] = 8'd194;
	sample_rom[204][4] = 8'd184;
	sample_rom[204][5] = 8'd177;
	sample_rom[204][6] = 8'd176;
	sample_rom[204][7] = 8'd180;
	sample_rom[204][8] = 8'd175;
	sample_rom[204][9] = 8'd165;
	sample_rom[204][10] = 8'd159;
	sample_rom[204][11] = 8'd156;
	sample_rom[204][12] = 8'd160;
	sample_rom[204][13] = 8'd162;
	sample_rom[204][14] = 8'd162;
	sample_rom[204][15] = 8'd157;
	sample_rom[204][16] = 8'd155;
	sample_rom[204][17] = 8'd155;
	sample_rom[204][18] = 8'd156;
	sample_rom[204][19] = 8'd150;
	sample_rom[204][20] = 8'd147;
	sample_rom[204][21] = 8'd145;
	sample_rom[204][22] = 8'd148;
	sample_rom[204][23] = 8'd151;
	sample_rom[204][24] = 8'd147;
	sample_rom[204][25] = 8'd145;
	sample_rom[204][26] = 8'd144;
	sample_rom[204][27] = 8'd145;
	sample_rom[204][28] = 8'd140;
	sample_rom[204][29] = 8'd145;
	sample_rom[204][30] = 8'd142;
	sample_rom[204][31] = 8'd138;
	sample_rom[204][32] = 8'd137;
	sample_rom[204][33] = 8'd140;
	sample_rom[204][34] = 8'd141;
	sample_rom[204][35] = 8'd136;
	sample_rom[204][36] = 8'd137;
	sample_rom[204][37] = 8'd133;
	sample_rom[204][38] = 8'd135;
	sample_rom[204][39] = 8'd131;
	sample_rom[204][40] = 8'd131;
	sample_rom[204][41] = 8'd128;
	sample_rom[204][42] = 8'd130;
	sample_rom[204][43] = 8'd131;
	sample_rom[204][44] = 8'd132;
	sample_rom[204][45] = 8'd133;
	sample_rom[204][46] = 8'd131;
	sample_rom[204][47] = 8'd134;
	sample_rom[204][48] = 8'd133;
	sample_rom[204][49] = 8'd131;
	sample_rom[204][50] = 8'd129;
	sample_rom[204][51] = 8'd128;
	sample_rom[204][52] = 8'd126;
	sample_rom[204][53] = 8'd128;
	sample_rom[204][54] = 8'd129;
	sample_rom[204][55] = 8'd129;
	sample_rom[204][56] = 8'd128;
	sample_rom[204][57] = 8'd125;
	sample_rom[204][58] = 8'd129;
	sample_rom[204][59] = 8'd128;
	sample_rom[204][60] = 8'd126;
	sample_rom[204][61] = 8'd130;
	sample_rom[204][62] = 8'd127;
	sample_rom[204][63] = 8'd127;
	sample_rom[205][0] = 8'd131;
	sample_rom[205][1] = 8'd210;
	sample_rom[205][2] = 8'd3;
	sample_rom[205][3] = 8'd10;
	sample_rom[205][4] = 8'd241;
	sample_rom[205][5] = 8'd224;
	sample_rom[205][6] = 8'd217;
	sample_rom[205][7] = 8'd216;
	sample_rom[205][8] = 8'd212;
	sample_rom[205][9] = 8'd200;
	sample_rom[205][10] = 8'd190;
	sample_rom[205][11] = 8'd188;
	sample_rom[205][12] = 8'd189;
	sample_rom[205][13] = 8'd186;
	sample_rom[205][14] = 8'd182;
	sample_rom[205][15] = 8'd177;
	sample_rom[205][16] = 8'd175;
	sample_rom[205][17] = 8'd174;
	sample_rom[205][18] = 8'd171;
	sample_rom[205][19] = 8'd171;
	sample_rom[205][20] = 8'd163;
	sample_rom[205][21] = 8'd161;
	sample_rom[205][22] = 8'd160;
	sample_rom[205][23] = 8'd162;
	sample_rom[205][24] = 8'd164;
	sample_rom[205][25] = 8'd153;
	sample_rom[205][26] = 8'd152;
	sample_rom[205][27] = 8'd147;
	sample_rom[205][28] = 8'd146;
	sample_rom[205][29] = 8'd153;
	sample_rom[205][30] = 8'd153;
	sample_rom[205][31] = 8'd148;
	sample_rom[205][32] = 8'd144;
	sample_rom[205][33] = 8'd144;
	sample_rom[205][34] = 8'd143;
	sample_rom[205][35] = 8'd145;
	sample_rom[205][36] = 8'd142;
	sample_rom[205][37] = 8'd138;
	sample_rom[205][38] = 8'd135;
	sample_rom[205][39] = 8'd132;
	sample_rom[205][40] = 8'd132;
	sample_rom[205][41] = 8'd130;
	sample_rom[205][42] = 8'd135;
	sample_rom[205][43] = 8'd136;
	sample_rom[205][44] = 8'd136;
	sample_rom[205][45] = 8'd134;
	sample_rom[205][46] = 8'd137;
	sample_rom[205][47] = 8'd138;
	sample_rom[205][48] = 8'd141;
	sample_rom[205][49] = 8'd141;
	sample_rom[205][50] = 8'd133;
	sample_rom[205][51] = 8'd129;
	sample_rom[205][52] = 8'd129;
	sample_rom[205][53] = 8'd127;
	sample_rom[205][54] = 8'd129;
	sample_rom[205][55] = 8'd127;
	sample_rom[205][56] = 8'd127;
	sample_rom[205][57] = 8'd125;
	sample_rom[205][58] = 8'd126;
	sample_rom[205][59] = 8'd127;
	sample_rom[205][60] = 8'd127;
	sample_rom[205][61] = 8'd126;
	sample_rom[205][62] = 8'd126;
	sample_rom[205][63] = 8'd128;
	sample_rom[206][0] = 8'd128;
	sample_rom[206][1] = 8'd170;
	sample_rom[206][2] = 8'd192;
	sample_rom[206][3] = 8'd191;
	sample_rom[206][4] = 8'd180;
	sample_rom[206][5] = 8'd173;
	sample_rom[206][6] = 8'd172;
	sample_rom[206][7] = 8'd175;
	sample_rom[206][8] = 8'd168;
	sample_rom[206][9] = 8'd159;
	sample_rom[206][10] = 8'd152;
	sample_rom[206][11] = 8'd149;
	sample_rom[206][12] = 8'd153;
	sample_rom[206][13] = 8'd154;
	sample_rom[206][14] = 8'd155;
	sample_rom[206][15] = 8'd149;
	sample_rom[206][16] = 8'd147;
	sample_rom[206][17] = 8'd147;
	sample_rom[206][18] = 8'd148;
	sample_rom[206][19] = 8'd143;
	sample_rom[206][20] = 8'd140;
	sample_rom[206][21] = 8'd139;
	sample_rom[206][22] = 8'd142;
	sample_rom[206][23] = 8'd145;
	sample_rom[206][24] = 8'd141;
	sample_rom[206][25] = 8'd140;
	sample_rom[206][26] = 8'd140;
	sample_rom[206][27] = 8'd141;
	sample_rom[206][28] = 8'd137;
	sample_rom[206][29] = 8'd141;
	sample_rom[206][30] = 8'd139;
	sample_rom[206][31] = 8'd135;
	sample_rom[206][32] = 8'd135;
	sample_rom[206][33] = 8'd138;
	sample_rom[206][34] = 8'd140;
	sample_rom[206][35] = 8'd134;
	sample_rom[206][36] = 8'd136;
	sample_rom[206][37] = 8'd132;
	sample_rom[206][38] = 8'd135;
	sample_rom[206][39] = 8'd130;
	sample_rom[206][40] = 8'd131;
	sample_rom[206][41] = 8'd129;
	sample_rom[206][42] = 8'd130;
	sample_rom[206][43] = 8'd131;
	sample_rom[206][44] = 8'd132;
	sample_rom[206][45] = 8'd133;
	sample_rom[206][46] = 8'd131;
	sample_rom[206][47] = 8'd134;
	sample_rom[206][48] = 8'd133;
	sample_rom[206][49] = 8'd132;
	sample_rom[206][50] = 8'd129;
	sample_rom[206][51] = 8'd127;
	sample_rom[206][52] = 8'd126;
	sample_rom[206][53] = 8'd127;
	sample_rom[206][54] = 8'd129;
	sample_rom[206][55] = 8'd128;
	sample_rom[206][56] = 8'd128;
	sample_rom[206][57] = 8'd125;
	sample_rom[206][58] = 8'd128;
	sample_rom[206][59] = 8'd127;
	sample_rom[206][60] = 8'd125;
	sample_rom[206][61] = 8'd130;
	sample_rom[206][62] = 8'd128;
	sample_rom[206][63] = 8'd126;
	sample_rom[207][0] = 8'd130;
	sample_rom[207][1] = 8'd212;
	sample_rom[207][2] = 8'd4;
	sample_rom[207][3] = 8'd2;
	sample_rom[207][4] = 8'd228;
	sample_rom[207][5] = 8'd216;
	sample_rom[207][6] = 8'd216;
	sample_rom[207][7] = 8'd220;
	sample_rom[207][8] = 8'd212;
	sample_rom[207][9] = 8'd190;
	sample_rom[207][10] = 8'd173;
	sample_rom[207][11] = 8'd172;
	sample_rom[207][12] = 8'd176;
	sample_rom[207][13] = 8'd178;
	sample_rom[207][14] = 8'd174;
	sample_rom[207][15] = 8'd167;
	sample_rom[207][16] = 8'd164;
	sample_rom[207][17] = 8'd167;
	sample_rom[207][18] = 8'd167;
	sample_rom[207][19] = 8'd164;
	sample_rom[207][20] = 8'd157;
	sample_rom[207][21] = 8'd151;
	sample_rom[207][22] = 8'd151;
	sample_rom[207][23] = 8'd158;
	sample_rom[207][24] = 8'd159;
	sample_rom[207][25] = 8'd150;
	sample_rom[207][26] = 8'd150;
	sample_rom[207][27] = 8'd147;
	sample_rom[207][28] = 8'd150;
	sample_rom[207][29] = 8'd150;
	sample_rom[207][30] = 8'd145;
	sample_rom[207][31] = 8'd142;
	sample_rom[207][32] = 8'd142;
	sample_rom[207][33] = 8'd147;
	sample_rom[207][34] = 8'd150;
	sample_rom[207][35] = 8'd148;
	sample_rom[207][36] = 8'd141;
	sample_rom[207][37] = 8'd138;
	sample_rom[207][38] = 8'd138;
	sample_rom[207][39] = 8'd133;
	sample_rom[207][40] = 8'd134;
	sample_rom[207][41] = 8'd128;
	sample_rom[207][42] = 8'd130;
	sample_rom[207][43] = 8'd133;
	sample_rom[207][44] = 8'd138;
	sample_rom[207][45] = 8'd139;
	sample_rom[207][46] = 8'd141;
	sample_rom[207][47] = 8'd135;
	sample_rom[207][48] = 8'd134;
	sample_rom[207][49] = 8'd138;
	sample_rom[207][50] = 8'd134;
	sample_rom[207][51] = 8'd127;
	sample_rom[207][52] = 8'd125;
	sample_rom[207][53] = 8'd124;
	sample_rom[207][54] = 8'd125;
	sample_rom[207][55] = 8'd126;
	sample_rom[207][56] = 8'd126;
	sample_rom[207][57] = 8'd122;
	sample_rom[207][58] = 8'd124;
	sample_rom[207][59] = 8'd126;
	sample_rom[207][60] = 8'd125;
	sample_rom[207][61] = 8'd125;
	sample_rom[207][62] = 8'd124;
	sample_rom[207][63] = 8'd129;
	sample_rom[208][0] = 8'd128;
	sample_rom[208][1] = 8'd170;
	sample_rom[208][2] = 8'd192;
	sample_rom[208][3] = 8'd191;
	sample_rom[208][4] = 8'd180;
	sample_rom[208][5] = 8'd173;
	sample_rom[208][6] = 8'd172;
	sample_rom[208][7] = 8'd175;
	sample_rom[208][8] = 8'd168;
	sample_rom[208][9] = 8'd159;
	sample_rom[208][10] = 8'd152;
	sample_rom[208][11] = 8'd149;
	sample_rom[208][12] = 8'd153;
	sample_rom[208][13] = 8'd154;
	sample_rom[208][14] = 8'd155;
	sample_rom[208][15] = 8'd149;
	sample_rom[208][16] = 8'd147;
	sample_rom[208][17] = 8'd147;
	sample_rom[208][18] = 8'd148;
	sample_rom[208][19] = 8'd143;
	sample_rom[208][20] = 8'd140;
	sample_rom[208][21] = 8'd139;
	sample_rom[208][22] = 8'd142;
	sample_rom[208][23] = 8'd145;
	sample_rom[208][24] = 8'd141;
	sample_rom[208][25] = 8'd140;
	sample_rom[208][26] = 8'd140;
	sample_rom[208][27] = 8'd141;
	sample_rom[208][28] = 8'd137;
	sample_rom[208][29] = 8'd141;
	sample_rom[208][30] = 8'd139;
	sample_rom[208][31] = 8'd135;
	sample_rom[208][32] = 8'd135;
	sample_rom[208][33] = 8'd138;
	sample_rom[208][34] = 8'd140;
	sample_rom[208][35] = 8'd134;
	sample_rom[208][36] = 8'd136;
	sample_rom[208][37] = 8'd132;
	sample_rom[208][38] = 8'd135;
	sample_rom[208][39] = 8'd130;
	sample_rom[208][40] = 8'd131;
	sample_rom[208][41] = 8'd129;
	sample_rom[208][42] = 8'd130;
	sample_rom[208][43] = 8'd131;
	sample_rom[208][44] = 8'd132;
	sample_rom[208][45] = 8'd133;
	sample_rom[208][46] = 8'd131;
	sample_rom[208][47] = 8'd134;
	sample_rom[208][48] = 8'd133;
	sample_rom[208][49] = 8'd132;
	sample_rom[208][50] = 8'd129;
	sample_rom[208][51] = 8'd127;
	sample_rom[208][52] = 8'd126;
	sample_rom[208][53] = 8'd127;
	sample_rom[208][54] = 8'd129;
	sample_rom[208][55] = 8'd128;
	sample_rom[208][56] = 8'd128;
	sample_rom[208][57] = 8'd125;
	sample_rom[208][58] = 8'd128;
	sample_rom[208][59] = 8'd127;
	sample_rom[208][60] = 8'd125;
	sample_rom[208][61] = 8'd130;
	sample_rom[208][62] = 8'd128;
	sample_rom[208][63] = 8'd126;
	sample_rom[209][0] = 8'd131;
	sample_rom[209][1] = 8'd139;
	sample_rom[209][2] = 8'd149;
	sample_rom[209][3] = 8'd158;
	sample_rom[209][4] = 8'd164;
	sample_rom[209][5] = 8'd173;
	sample_rom[209][6] = 8'd179;
	sample_rom[209][7] = 8'd186;
	sample_rom[209][8] = 8'd191;
	sample_rom[209][9] = 8'd195;
	sample_rom[209][10] = 8'd200;
	sample_rom[209][11] = 8'd203;
	sample_rom[209][12] = 8'd205;
	sample_rom[209][13] = 8'd207;
	sample_rom[209][14] = 8'd208;
	sample_rom[209][15] = 8'd208;
	sample_rom[209][16] = 8'd207;
	sample_rom[209][17] = 8'd204;
	sample_rom[209][18] = 8'd202;
	sample_rom[209][19] = 8'd199;
	sample_rom[209][20] = 8'd194;
	sample_rom[209][21] = 8'd191;
	sample_rom[209][22] = 8'd185;
	sample_rom[209][23] = 8'd180;
	sample_rom[209][24] = 8'd175;
	sample_rom[209][25] = 8'd168;
	sample_rom[209][26] = 8'd163;
	sample_rom[209][27] = 8'd159;
	sample_rom[209][28] = 8'd153;
	sample_rom[209][29] = 8'd149;
	sample_rom[209][30] = 8'd144;
	sample_rom[209][31] = 8'd139;
	sample_rom[209][32] = 8'd135;
	sample_rom[209][33] = 8'd132;
	sample_rom[209][34] = 8'd128;
	sample_rom[209][35] = 8'd126;
	sample_rom[209][36] = 8'd124;
	sample_rom[209][37] = 8'd122;
	sample_rom[209][38] = 8'd120;
	sample_rom[209][39] = 8'd120;
	sample_rom[209][40] = 8'd119;
	sample_rom[209][41] = 8'd120;
	sample_rom[209][42] = 8'd121;
	sample_rom[209][43] = 8'd122;
	sample_rom[209][44] = 8'd122;
	sample_rom[209][45] = 8'd124;
	sample_rom[209][46] = 8'd125;
	sample_rom[209][47] = 8'd126;
	sample_rom[209][48] = 8'd127;
	sample_rom[209][49] = 8'd130;
	sample_rom[209][50] = 8'd130;
	sample_rom[209][51] = 8'd131;
	sample_rom[209][52] = 8'd132;
	sample_rom[209][53] = 8'd133;
	sample_rom[209][54] = 8'd134;
	sample_rom[209][55] = 8'd134;
	sample_rom[209][56] = 8'd135;
	sample_rom[209][57] = 8'd134;
	sample_rom[209][58] = 8'd134;
	sample_rom[209][59] = 8'd133;
	sample_rom[209][60] = 8'd133;
	sample_rom[209][61] = 8'd131;
	sample_rom[209][62] = 8'd129;
	sample_rom[209][63] = 8'd129;
	sample_rom[210][0] = 8'd132;
	sample_rom[210][1] = 8'd145;
	sample_rom[210][2] = 8'd157;
	sample_rom[210][3] = 8'd168;
	sample_rom[210][4] = 8'd178;
	sample_rom[210][5] = 8'd189;
	sample_rom[210][6] = 8'd198;
	sample_rom[210][7] = 8'd207;
	sample_rom[210][8] = 8'd215;
	sample_rom[210][9] = 8'd222;
	sample_rom[210][10] = 8'd226;
	sample_rom[210][11] = 8'd231;
	sample_rom[210][12] = 8'd234;
	sample_rom[210][13] = 8'd235;
	sample_rom[210][14] = 8'd235;
	sample_rom[210][15] = 8'd235;
	sample_rom[210][16] = 8'd233;
	sample_rom[210][17] = 8'd230;
	sample_rom[210][18] = 8'd226;
	sample_rom[210][19] = 8'd222;
	sample_rom[210][20] = 8'd217;
	sample_rom[210][21] = 8'd211;
	sample_rom[210][22] = 8'd205;
	sample_rom[210][23] = 8'd198;
	sample_rom[210][24] = 8'd191;
	sample_rom[210][25] = 8'd185;
	sample_rom[210][26] = 8'd178;
	sample_rom[210][27] = 8'd172;
	sample_rom[210][28] = 8'd166;
	sample_rom[210][29] = 8'd161;
	sample_rom[210][30] = 8'd158;
	sample_rom[210][31] = 8'd154;
	sample_rom[210][32] = 8'd150;
	sample_rom[210][33] = 8'd149;
	sample_rom[210][34] = 8'd147;
	sample_rom[210][35] = 8'd146;
	sample_rom[210][36] = 8'd147;
	sample_rom[210][37] = 8'd147;
	sample_rom[210][38] = 8'd149;
	sample_rom[210][39] = 8'd151;
	sample_rom[210][40] = 8'd154;
	sample_rom[210][41] = 8'd156;
	sample_rom[210][42] = 8'd160;
	sample_rom[210][43] = 8'd162;
	sample_rom[210][44] = 8'd166;
	sample_rom[210][45] = 8'd169;
	sample_rom[210][46] = 8'd173;
	sample_rom[210][47] = 8'd175;
	sample_rom[210][48] = 8'd178;
	sample_rom[210][49] = 8'd179;
	sample_rom[210][50] = 8'd180;
	sample_rom[210][51] = 8'd182;
	sample_rom[210][52] = 8'd181;
	sample_rom[210][53] = 8'd180;
	sample_rom[210][54] = 8'd177;
	sample_rom[210][55] = 8'd175;
	sample_rom[210][56] = 8'd172;
	sample_rom[210][57] = 8'd168;
	sample_rom[210][58] = 8'd163;
	sample_rom[210][59] = 8'd160;
	sample_rom[210][60] = 8'd153;
	sample_rom[210][61] = 8'd148;
	sample_rom[210][62] = 8'd140;
	sample_rom[210][63] = 8'd134;
	sample_rom[211][0] = 8'd132;
	sample_rom[211][1] = 8'd142;
	sample_rom[211][2] = 8'd154;
	sample_rom[211][3] = 8'd164;
	sample_rom[211][4] = 8'd173;
	sample_rom[211][5] = 8'd183;
	sample_rom[211][6] = 8'd191;
	sample_rom[211][7] = 8'd199;
	sample_rom[211][8] = 8'd205;
	sample_rom[211][9] = 8'd211;
	sample_rom[211][10] = 8'd217;
	sample_rom[211][11] = 8'd222;
	sample_rom[211][12] = 8'd223;
	sample_rom[211][13] = 8'd225;
	sample_rom[211][14] = 8'd228;
	sample_rom[211][15] = 8'd229;
	sample_rom[211][16] = 8'd229;
	sample_rom[211][17] = 8'd228;
	sample_rom[211][18] = 8'd228;
	sample_rom[211][19] = 8'd227;
	sample_rom[211][20] = 8'd224;
	sample_rom[211][21] = 8'd224;
	sample_rom[211][22] = 8'd223;
	sample_rom[211][23] = 8'd222;
	sample_rom[211][24] = 8'd220;
	sample_rom[211][25] = 8'd219;
	sample_rom[211][26] = 8'd218;
	sample_rom[211][27] = 8'd219;
	sample_rom[211][28] = 8'd219;
	sample_rom[211][29] = 8'd219;
	sample_rom[211][30] = 8'd220;
	sample_rom[211][31] = 8'd221;
	sample_rom[211][32] = 8'd222;
	sample_rom[211][33] = 8'd224;
	sample_rom[211][34] = 8'd224;
	sample_rom[211][35] = 8'd227;
	sample_rom[211][36] = 8'd229;
	sample_rom[211][37] = 8'd230;
	sample_rom[211][38] = 8'd231;
	sample_rom[211][39] = 8'd233;
	sample_rom[211][40] = 8'd234;
	sample_rom[211][41] = 8'd235;
	sample_rom[211][42] = 8'd235;
	sample_rom[211][43] = 8'd235;
	sample_rom[211][44] = 8'd235;
	sample_rom[211][45] = 8'd233;
	sample_rom[211][46] = 8'd231;
	sample_rom[211][47] = 8'd228;
	sample_rom[211][48] = 8'd226;
	sample_rom[211][49] = 8'd223;
	sample_rom[211][50] = 8'd218;
	sample_rom[211][51] = 8'd213;
	sample_rom[211][52] = 8'd208;
	sample_rom[211][53] = 8'd203;
	sample_rom[211][54] = 8'd197;
	sample_rom[211][55] = 8'd190;
	sample_rom[211][56] = 8'd184;
	sample_rom[211][57] = 8'd177;
	sample_rom[211][58] = 8'd170;
	sample_rom[211][59] = 8'd163;
	sample_rom[211][60] = 8'd157;
	sample_rom[211][61] = 8'd149;
	sample_rom[211][62] = 8'd139;
	sample_rom[211][63] = 8'd133;
	sample_rom[212][0] = 8'd132;
	sample_rom[212][1] = 8'd150;
	sample_rom[212][2] = 8'd164;
	sample_rom[212][3] = 8'd179;
	sample_rom[212][4] = 8'd194;
	sample_rom[212][5] = 8'd206;
	sample_rom[212][6] = 8'd216;
	sample_rom[212][7] = 8'd224;
	sample_rom[212][8] = 8'd230;
	sample_rom[212][9] = 8'd233;
	sample_rom[212][10] = 8'd234;
	sample_rom[212][11] = 8'd231;
	sample_rom[212][12] = 8'd227;
	sample_rom[212][13] = 8'd222;
	sample_rom[212][14] = 8'd214;
	sample_rom[212][15] = 8'd204;
	sample_rom[212][16] = 8'd194;
	sample_rom[212][17] = 8'd183;
	sample_rom[212][18] = 8'd172;
	sample_rom[212][19] = 8'd162;
	sample_rom[212][20] = 8'd154;
	sample_rom[212][21] = 8'd145;
	sample_rom[212][22] = 8'd137;
	sample_rom[212][23] = 8'd131;
	sample_rom[212][24] = 8'd126;
	sample_rom[212][25] = 8'd126;
	sample_rom[212][26] = 8'd125;
	sample_rom[212][27] = 8'd127;
	sample_rom[212][28] = 8'd131;
	sample_rom[212][29] = 8'd137;
	sample_rom[212][30] = 8'd145;
	sample_rom[212][31] = 8'd153;
	sample_rom[212][32] = 8'd160;
	sample_rom[212][33] = 8'd171;
	sample_rom[212][34] = 8'd179;
	sample_rom[212][35] = 8'd189;
	sample_rom[212][36] = 8'd198;
	sample_rom[212][37] = 8'd205;
	sample_rom[212][38] = 8'd213;
	sample_rom[212][39] = 8'd217;
	sample_rom[212][40] = 8'd222;
	sample_rom[212][41] = 8'd223;
	sample_rom[212][42] = 8'd224;
	sample_rom[212][43] = 8'd222;
	sample_rom[212][44] = 8'd219;
	sample_rom[212][45] = 8'd215;
	sample_rom[212][46] = 8'd208;
	sample_rom[212][47] = 8'd201;
	sample_rom[212][48] = 8'd193;
	sample_rom[212][49] = 8'd185;
	sample_rom[212][50] = 8'd175;
	sample_rom[212][51] = 8'd167;
	sample_rom[212][52] = 8'd159;
	sample_rom[212][53] = 8'd152;
	sample_rom[212][54] = 8'd145;
	sample_rom[212][55] = 8'd138;
	sample_rom[212][56] = 8'd132;
	sample_rom[212][57] = 8'd129;
	sample_rom[212][58] = 8'd126;
	sample_rom[212][59] = 8'd124;
	sample_rom[212][60] = 8'd123;
	sample_rom[212][61] = 8'd124;
	sample_rom[212][62] = 8'd125;
	sample_rom[212][63] = 8'd126;
	sample_rom[213][0] = 8'd132;
	sample_rom[213][1] = 8'd150;
	sample_rom[213][2] = 8'd168;
	sample_rom[213][3] = 8'd185;
	sample_rom[213][4] = 8'd201;
	sample_rom[213][5] = 8'd215;
	sample_rom[213][6] = 8'd226;
	sample_rom[213][7] = 8'd235;
	sample_rom[213][8] = 8'd243;
	sample_rom[213][9] = 8'd248;
	sample_rom[213][10] = 8'd251;
	sample_rom[213][11] = 8'd251;
	sample_rom[213][12] = 8'd248;
	sample_rom[213][13] = 8'd242;
	sample_rom[213][14] = 8'd235;
	sample_rom[213][15] = 8'd226;
	sample_rom[213][16] = 8'd216;
	sample_rom[213][17] = 8'd204;
	sample_rom[213][18] = 8'd191;
	sample_rom[213][19] = 8'd177;
	sample_rom[213][20] = 8'd164;
	sample_rom[213][21] = 8'd152;
	sample_rom[213][22] = 8'd138;
	sample_rom[213][23] = 8'd128;
	sample_rom[213][24] = 8'd116;
	sample_rom[213][25] = 8'd108;
	sample_rom[213][26] = 8'd100;
	sample_rom[213][27] = 8'd97;
	sample_rom[213][28] = 8'd93;
	sample_rom[213][29] = 8'd91;
	sample_rom[213][30] = 8'd92;
	sample_rom[213][31] = 8'd94;
	sample_rom[213][32] = 8'd98;
	sample_rom[213][33] = 8'd103;
	sample_rom[213][34] = 8'd109;
	sample_rom[213][35] = 8'd118;
	sample_rom[213][36] = 8'd127;
	sample_rom[213][37] = 8'd137;
	sample_rom[213][38] = 8'd146;
	sample_rom[213][39] = 8'd156;
	sample_rom[213][40] = 8'd166;
	sample_rom[213][41] = 8'd175;
	sample_rom[213][42] = 8'd185;
	sample_rom[213][43] = 8'd193;
	sample_rom[213][44] = 8'd201;
	sample_rom[213][45] = 8'd207;
	sample_rom[213][46] = 8'd211;
	sample_rom[213][47] = 8'd215;
	sample_rom[213][48] = 8'd217;
	sample_rom[213][49] = 8'd218;
	sample_rom[213][50] = 8'd217;
	sample_rom[213][51] = 8'd216;
	sample_rom[213][52] = 8'd214;
	sample_rom[213][53] = 8'd210;
	sample_rom[213][54] = 8'd205;
	sample_rom[213][55] = 8'd199;
	sample_rom[213][56] = 8'd193;
	sample_rom[213][57] = 8'd186;
	sample_rom[213][58] = 8'd178;
	sample_rom[213][59] = 8'd171;
	sample_rom[213][60] = 8'd162;
	sample_rom[213][61] = 8'd153;
	sample_rom[213][62] = 8'd143;
	sample_rom[213][63] = 8'd135;
	sample_rom[214][0] = 8'd132;
	sample_rom[214][1] = 8'd153;
	sample_rom[214][2] = 8'd173;
	sample_rom[214][3] = 8'd191;
	sample_rom[214][4] = 8'd205;
	sample_rom[214][5] = 8'd217;
	sample_rom[214][6] = 8'd224;
	sample_rom[214][7] = 8'd227;
	sample_rom[214][8] = 8'd227;
	sample_rom[214][9] = 8'd223;
	sample_rom[214][10] = 8'd215;
	sample_rom[214][11] = 8'd203;
	sample_rom[214][12] = 8'd191;
	sample_rom[214][13] = 8'd175;
	sample_rom[214][14] = 8'd161;
	sample_rom[214][15] = 8'd146;
	sample_rom[214][16] = 8'd133;
	sample_rom[214][17] = 8'd122;
	sample_rom[214][18] = 8'd115;
	sample_rom[214][19] = 8'd110;
	sample_rom[214][20] = 8'd111;
	sample_rom[214][21] = 8'd115;
	sample_rom[214][22] = 8'd121;
	sample_rom[214][23] = 8'd131;
	sample_rom[214][24] = 8'd143;
	sample_rom[214][25] = 8'd159;
	sample_rom[214][26] = 8'd173;
	sample_rom[214][27] = 8'd190;
	sample_rom[214][28] = 8'd206;
	sample_rom[214][29] = 8'd219;
	sample_rom[214][30] = 8'd230;
	sample_rom[214][31] = 8'd240;
	sample_rom[214][32] = 8'd247;
	sample_rom[214][33] = 8'd248;
	sample_rom[214][34] = 8'd248;
	sample_rom[214][35] = 8'd243;
	sample_rom[214][36] = 8'd235;
	sample_rom[214][37] = 8'd225;
	sample_rom[214][38] = 8'd214;
	sample_rom[214][39] = 8'd199;
	sample_rom[214][40] = 8'd187;
	sample_rom[214][41] = 8'd173;
	sample_rom[214][42] = 8'd161;
	sample_rom[214][43] = 8'd151;
	sample_rom[214][44] = 8'd142;
	sample_rom[214][45] = 8'd135;
	sample_rom[214][46] = 8'd132;
	sample_rom[214][47] = 8'd131;
	sample_rom[214][48] = 8'd133;
	sample_rom[214][49] = 8'd137;
	sample_rom[214][50] = 8'd142;
	sample_rom[214][51] = 8'd150;
	sample_rom[214][52] = 8'd157;
	sample_rom[214][53] = 8'd164;
	sample_rom[214][54] = 8'd170;
	sample_rom[214][55] = 8'd176;
	sample_rom[214][56] = 8'd178;
	sample_rom[214][57] = 8'd179;
	sample_rom[214][58] = 8'd177;
	sample_rom[214][59] = 8'd174;
	sample_rom[214][60] = 8'd168;
	sample_rom[214][61] = 8'd159;
	sample_rom[214][62] = 8'd149;
	sample_rom[214][63] = 8'd138;
	sample_rom[215][0] = 8'd130;
	sample_rom[215][1] = 8'd149;
	sample_rom[215][2] = 8'd166;
	sample_rom[215][3] = 8'd179;
	sample_rom[215][4] = 8'd192;
	sample_rom[215][5] = 8'd203;
	sample_rom[215][6] = 8'd209;
	sample_rom[215][7] = 8'd216;
	sample_rom[215][8] = 8'd217;
	sample_rom[215][9] = 8'd216;
	sample_rom[215][10] = 8'd214;
	sample_rom[215][11] = 8'd209;
	sample_rom[215][12] = 8'd203;
	sample_rom[215][13] = 8'd198;
	sample_rom[215][14] = 8'd192;
	sample_rom[215][15] = 8'd187;
	sample_rom[215][16] = 8'd183;
	sample_rom[215][17] = 8'd177;
	sample_rom[215][18] = 8'd177;
	sample_rom[215][19] = 8'd179;
	sample_rom[215][20] = 8'd179;
	sample_rom[215][21] = 8'd183;
	sample_rom[215][22] = 8'd188;
	sample_rom[215][23] = 8'd194;
	sample_rom[215][24] = 8'd199;
	sample_rom[215][25] = 8'd206;
	sample_rom[215][26] = 8'd211;
	sample_rom[215][27] = 8'd217;
	sample_rom[215][28] = 8'd220;
	sample_rom[215][29] = 8'd223;
	sample_rom[215][30] = 8'd224;
	sample_rom[215][31] = 8'd224;
	sample_rom[215][32] = 8'd223;
	sample_rom[215][33] = 8'd223;
	sample_rom[215][34] = 8'd219;
	sample_rom[215][35] = 8'd217;
	sample_rom[215][36] = 8'd213;
	sample_rom[215][37] = 8'd208;
	sample_rom[215][38] = 8'd204;
	sample_rom[215][39] = 8'd201;
	sample_rom[215][40] = 8'd199;
	sample_rom[215][41] = 8'd195;
	sample_rom[215][42] = 8'd193;
	sample_rom[215][43] = 8'd189;
	sample_rom[215][44] = 8'd187;
	sample_rom[215][45] = 8'd184;
	sample_rom[215][46] = 8'd179;
	sample_rom[215][47] = 8'd176;
	sample_rom[215][48] = 8'd171;
	sample_rom[215][49] = 8'd167;
	sample_rom[215][50] = 8'd160;
	sample_rom[215][51] = 8'd154;
	sample_rom[215][52] = 8'd149;
	sample_rom[215][53] = 8'd143;
	sample_rom[215][54] = 8'd137;
	sample_rom[215][55] = 8'd132;
	sample_rom[215][56] = 8'd126;
	sample_rom[215][57] = 8'd123;
	sample_rom[215][58] = 8'd121;
	sample_rom[215][59] = 8'd120;
	sample_rom[215][60] = 8'd121;
	sample_rom[215][61] = 8'd121;
	sample_rom[215][62] = 8'd122;
	sample_rom[215][63] = 8'd124;
	sample_rom[216][0] = 8'd131;
	sample_rom[216][1] = 8'd154;
	sample_rom[216][2] = 8'd174;
	sample_rom[216][3] = 8'd192;
	sample_rom[216][4] = 8'd208;
	sample_rom[216][5] = 8'd219;
	sample_rom[216][6] = 8'd227;
	sample_rom[216][7] = 8'd230;
	sample_rom[216][8] = 8'd228;
	sample_rom[216][9] = 8'd223;
	sample_rom[216][10] = 8'd218;
	sample_rom[216][11] = 8'd208;
	sample_rom[216][12] = 8'd198;
	sample_rom[216][13] = 8'd188;
	sample_rom[216][14] = 8'd178;
	sample_rom[216][15] = 8'd171;
	sample_rom[216][16] = 8'd167;
	sample_rom[216][17] = 8'd161;
	sample_rom[216][18] = 8'd164;
	sample_rom[216][19] = 8'd164;
	sample_rom[216][20] = 8'd169;
	sample_rom[216][21] = 8'd177;
	sample_rom[216][22] = 8'd183;
	sample_rom[216][23] = 8'd191;
	sample_rom[216][24] = 8'd196;
	sample_rom[216][25] = 8'd202;
	sample_rom[216][26] = 8'd205;
	sample_rom[216][27] = 8'd204;
	sample_rom[216][28] = 8'd203;
	sample_rom[216][29] = 8'd198;
	sample_rom[216][30] = 8'd192;
	sample_rom[216][31] = 8'd184;
	sample_rom[216][32] = 8'd172;
	sample_rom[216][33] = 8'd162;
	sample_rom[216][34] = 8'd152;
	sample_rom[216][35] = 8'd143;
	sample_rom[216][36] = 8'd135;
	sample_rom[216][37] = 8'd129;
	sample_rom[216][38] = 8'd124;
	sample_rom[216][39] = 8'd122;
	sample_rom[216][40] = 8'd123;
	sample_rom[216][41] = 8'd124;
	sample_rom[216][42] = 8'd126;
	sample_rom[216][43] = 8'd129;
	sample_rom[216][44] = 8'd131;
	sample_rom[216][45] = 8'd133;
	sample_rom[216][46] = 8'd134;
	sample_rom[216][47] = 8'd134;
	sample_rom[216][48] = 8'd130;
	sample_rom[216][49] = 8'd126;
	sample_rom[216][50] = 8'd120;
	sample_rom[216][51] = 8'd111;
	sample_rom[216][52] = 8'd102;
	sample_rom[216][53] = 8'd93;
	sample_rom[216][54] = 8'd86;
	sample_rom[216][55] = 8'd78;
	sample_rom[216][56] = 8'd72;
	sample_rom[216][57] = 8'd70;
	sample_rom[216][58] = 8'd70;
	sample_rom[216][59] = 8'd75;
	sample_rom[216][60] = 8'd82;
	sample_rom[216][61] = 8'd92;
	sample_rom[216][62] = 8'd103;
	sample_rom[216][63] = 8'd115;
	sample_rom[217][0] = 8'd131;
	sample_rom[217][1] = 8'd166;
	sample_rom[217][2] = 8'd197;
	sample_rom[217][3] = 8'd222;
	sample_rom[217][4] = 8'd238;
	sample_rom[217][5] = 8'd250;
	sample_rom[217][6] = 8'd248;
	sample_rom[217][7] = 8'd241;
	sample_rom[217][8] = 8'd226;
	sample_rom[217][9] = 8'd206;
	sample_rom[217][10] = 8'd185;
	sample_rom[217][11] = 8'd162;
	sample_rom[217][12] = 8'd144;
	sample_rom[217][13] = 8'd128;
	sample_rom[217][14] = 8'd118;
	sample_rom[217][15] = 8'd116;
	sample_rom[217][16] = 8'd116;
	sample_rom[217][17] = 8'd126;
	sample_rom[217][18] = 8'd138;
	sample_rom[217][19] = 8'd153;
	sample_rom[217][20] = 8'd167;
	sample_rom[217][21] = 8'd180;
	sample_rom[217][22] = 8'd192;
	sample_rom[217][23] = 8'd198;
	sample_rom[217][24] = 8'd200;
	sample_rom[217][25] = 8'd197;
	sample_rom[217][26] = 8'd190;
	sample_rom[217][27] = 8'd180;
	sample_rom[217][28] = 8'd167;
	sample_rom[217][29] = 8'd155;
	sample_rom[217][30] = 8'd142;
	sample_rom[217][31] = 8'd132;
	sample_rom[217][32] = 8'd123;
	sample_rom[217][33] = 8'd117;
	sample_rom[217][34] = 8'd112;
	sample_rom[217][35] = 8'd112;
	sample_rom[217][36] = 8'd111;
	sample_rom[217][37] = 8'd111;
	sample_rom[217][38] = 8'd111;
	sample_rom[217][39] = 8'd106;
	sample_rom[217][40] = 8'd102;
	sample_rom[217][41] = 8'd95;
	sample_rom[217][42] = 8'd86;
	sample_rom[217][43] = 8'd74;
	sample_rom[217][44] = 8'd62;
	sample_rom[217][45] = 8'd51;
	sample_rom[217][46] = 8'd37;
	sample_rom[217][47] = 8'd31;
	sample_rom[217][48] = 8'd26;
	sample_rom[217][49] = 8'd29;
	sample_rom[217][50] = 8'd34;
	sample_rom[217][51] = 8'd43;
	sample_rom[217][52] = 8'd60;
	sample_rom[217][53] = 8'd77;
	sample_rom[217][54] = 8'd96;
	sample_rom[217][55] = 8'd113;
	sample_rom[217][56] = 8'd133;
	sample_rom[217][57] = 8'd148;
	sample_rom[217][58] = 8'd158;
	sample_rom[217][59] = 8'd164;
	sample_rom[217][60] = 8'd164;
	sample_rom[217][61] = 8'd160;
	sample_rom[217][62] = 8'd152;
	sample_rom[217][63] = 8'd142;
	sample_rom[218][0] = 8'd131;
	sample_rom[218][1] = 8'd164;
	sample_rom[218][2] = 8'd196;
	sample_rom[218][3] = 8'd217;
	sample_rom[218][4] = 8'd228;
	sample_rom[218][5] = 8'd233;
	sample_rom[218][6] = 8'd224;
	sample_rom[218][7] = 8'd211;
	sample_rom[218][8] = 8'd187;
	sample_rom[218][9] = 8'd165;
	sample_rom[218][10] = 8'd143;
	sample_rom[218][11] = 8'd124;
	sample_rom[218][12] = 8'd113;
	sample_rom[218][13] = 8'd109;
	sample_rom[218][14] = 8'd114;
	sample_rom[218][15] = 8'd127;
	sample_rom[218][16] = 8'd145;
	sample_rom[218][17] = 8'd165;
	sample_rom[218][18] = 8'd186;
	sample_rom[218][19] = 8'd203;
	sample_rom[218][20] = 8'd214;
	sample_rom[218][21] = 8'd218;
	sample_rom[218][22] = 8'd215;
	sample_rom[218][23] = 8'd206;
	sample_rom[218][24] = 8'd190;
	sample_rom[218][25] = 8'd171;
	sample_rom[218][26] = 8'd150;
	sample_rom[218][27] = 8'd132;
	sample_rom[218][28] = 8'd117;
	sample_rom[218][29] = 8'd108;
	sample_rom[218][30] = 8'd102;
	sample_rom[218][31] = 8'd100;
	sample_rom[218][32] = 8'd104;
	sample_rom[218][33] = 8'd110;
	sample_rom[218][34] = 8'd116;
	sample_rom[218][35] = 8'd120;
	sample_rom[218][36] = 8'd121;
	sample_rom[218][37] = 8'd119;
	sample_rom[218][38] = 8'd111;
	sample_rom[218][39] = 8'd103;
	sample_rom[218][40] = 8'd92;
	sample_rom[218][41] = 8'd84;
	sample_rom[218][42] = 8'd73;
	sample_rom[218][43] = 8'd67;
	sample_rom[218][44] = 8'd65;
	sample_rom[218][45] = 8'd69;
	sample_rom[218][46] = 8'd76;
	sample_rom[218][47] = 8'd86;
	sample_rom[218][48] = 8'd97;
	sample_rom[218][49] = 8'd110;
	sample_rom[218][50] = 8'd119;
	sample_rom[218][51] = 8'd126;
	sample_rom[218][52] = 8'd128;
	sample_rom[218][53] = 8'd123;
	sample_rom[218][54] = 8'd114;
	sample_rom[218][55] = 8'd104;
	sample_rom[218][56] = 8'd91;
	sample_rom[218][57] = 8'd80;
	sample_rom[218][58] = 8'd71;
	sample_rom[218][59] = 8'd68;
	sample_rom[218][60] = 8'd70;
	sample_rom[218][61] = 8'd80;
	sample_rom[218][62] = 8'd94;
	sample_rom[218][63] = 8'd110;
	sample_rom[219][0] = 8'd130;
	sample_rom[219][1] = 8'd163;
	sample_rom[219][2] = 8'd191;
	sample_rom[219][3] = 8'd212;
	sample_rom[219][4] = 8'd225;
	sample_rom[219][5] = 8'd230;
	sample_rom[219][6] = 8'd225;
	sample_rom[219][7] = 8'd215;
	sample_rom[219][8] = 8'd199;
	sample_rom[219][9] = 8'd182;
	sample_rom[219][10] = 8'd165;
	sample_rom[219][11] = 8'd154;
	sample_rom[219][12] = 8'd145;
	sample_rom[219][13] = 8'd143;
	sample_rom[219][14] = 8'd144;
	sample_rom[219][15] = 8'd151;
	sample_rom[219][16] = 8'd159;
	sample_rom[219][17] = 8'd163;
	sample_rom[219][18] = 8'd166;
	sample_rom[219][19] = 8'd168;
	sample_rom[219][20] = 8'd166;
	sample_rom[219][21] = 8'd160;
	sample_rom[219][22] = 8'd151;
	sample_rom[219][23] = 8'd142;
	sample_rom[219][24] = 8'd132;
	sample_rom[219][25] = 8'd122;
	sample_rom[219][26] = 8'd116;
	sample_rom[219][27] = 8'd111;
	sample_rom[219][28] = 8'd108;
	sample_rom[219][29] = 8'd105;
	sample_rom[219][30] = 8'd103;
	sample_rom[219][31] = 8'd99;
	sample_rom[219][32] = 8'd93;
	sample_rom[219][33] = 8'd86;
	sample_rom[219][34] = 8'd76;
	sample_rom[219][35] = 8'd69;
	sample_rom[219][36] = 8'd60;
	sample_rom[219][37] = 8'd54;
	sample_rom[219][38] = 8'd54;
	sample_rom[219][39] = 8'd58;
	sample_rom[219][40] = 8'd68;
	sample_rom[219][41] = 8'd85;
	sample_rom[219][42] = 8'd102;
	sample_rom[219][43] = 8'd123;
	sample_rom[219][44] = 8'd143;
	sample_rom[219][45] = 8'd159;
	sample_rom[219][46] = 8'd173;
	sample_rom[219][47] = 8'd178;
	sample_rom[219][48] = 8'd180;
	sample_rom[219][49] = 8'd179;
	sample_rom[219][50] = 8'd170;
	sample_rom[219][51] = 8'd162;
	sample_rom[219][52] = 8'd154;
	sample_rom[219][53] = 8'd145;
	sample_rom[219][54] = 8'd139;
	sample_rom[219][55] = 8'd135;
	sample_rom[219][56] = 8'd135;
	sample_rom[219][57] = 8'd136;
	sample_rom[219][58] = 8'd138;
	sample_rom[219][59] = 8'd140;
	sample_rom[219][60] = 8'd140;
	sample_rom[219][61] = 8'd139;
	sample_rom[219][62] = 8'd137;
	sample_rom[219][63] = 8'd133;
	sample_rom[220][0] = 8'd132;
	sample_rom[220][1] = 8'd176;
	sample_rom[220][2] = 8'd213;
	sample_rom[220][3] = 8'd239;
	sample_rom[220][4] = 8'd250;
	sample_rom[220][5] = 8'd250;
	sample_rom[220][6] = 8'd236;
	sample_rom[220][7] = 8'd218;
	sample_rom[220][8] = 8'd196;
	sample_rom[220][9] = 8'd178;
	sample_rom[220][10] = 8'd172;
	sample_rom[220][11] = 8'd172;
	sample_rom[220][12] = 8'd181;
	sample_rom[220][13] = 8'd197;
	sample_rom[220][14] = 8'd213;
	sample_rom[220][15] = 8'd225;
	sample_rom[220][16] = 8'd233;
	sample_rom[220][17] = 8'd231;
	sample_rom[220][18] = 8'd221;
	sample_rom[220][19] = 8'd204;
	sample_rom[220][20] = 8'd182;
	sample_rom[220][21] = 8'd160;
	sample_rom[220][22] = 8'd138;
	sample_rom[220][23] = 8'd122;
	sample_rom[220][24] = 8'd111;
	sample_rom[220][25] = 8'd101;
	sample_rom[220][26] = 8'd98;
	sample_rom[220][27] = 8'd94;
	sample_rom[220][28] = 8'd88;
	sample_rom[220][29] = 8'd81;
	sample_rom[220][30] = 8'd70;
	sample_rom[220][31] = 8'd57;
	sample_rom[220][32] = 8'd43;
	sample_rom[220][33] = 8'd34;
	sample_rom[220][34] = 8'd29;
	sample_rom[220][35] = 8'd33;
	sample_rom[220][36] = 8'd42;
	sample_rom[220][37] = 8'd55;
	sample_rom[220][38] = 8'd73;
	sample_rom[220][39] = 8'd91;
	sample_rom[220][40] = 8'd109;
	sample_rom[220][41] = 8'd118;
	sample_rom[220][42] = 8'd127;
	sample_rom[220][43] = 8'd129;
	sample_rom[220][44] = 8'd128;
	sample_rom[220][45] = 8'd123;
	sample_rom[220][46] = 8'd119;
	sample_rom[220][47] = 8'd117;
	sample_rom[220][48] = 8'd120;
	sample_rom[220][49] = 8'd130;
	sample_rom[220][50] = 8'd141;
	sample_rom[220][51] = 8'd156;
	sample_rom[220][52] = 8'd169;
	sample_rom[220][53] = 8'd182;
	sample_rom[220][54] = 8'd189;
	sample_rom[220][55] = 8'd193;
	sample_rom[220][56] = 8'd193;
	sample_rom[220][57] = 8'd183;
	sample_rom[220][58] = 8'd176;
	sample_rom[220][59] = 8'd162;
	sample_rom[220][60] = 8'd152;
	sample_rom[220][61] = 8'd143;
	sample_rom[220][62] = 8'd136;
	sample_rom[220][63] = 8'd133;
	sample_rom[221][0] = 8'd131;
	sample_rom[221][1] = 8'd179;
	sample_rom[221][2] = 8'd216;
	sample_rom[221][3] = 8'd237;
	sample_rom[221][4] = 8'd241;
	sample_rom[221][5] = 8'd226;
	sample_rom[221][6] = 8'd204;
	sample_rom[221][7] = 8'd179;
	sample_rom[221][8] = 8'd161;
	sample_rom[221][9] = 8'd156;
	sample_rom[221][10] = 8'd162;
	sample_rom[221][11] = 8'd180;
	sample_rom[221][12] = 8'd207;
	sample_rom[221][13] = 8'd230;
	sample_rom[221][14] = 8'd246;
	sample_rom[221][15] = 8'd251;
	sample_rom[221][16] = 8'd241;
	sample_rom[221][17] = 8'd222;
	sample_rom[221][18] = 8'd198;
	sample_rom[221][19] = 8'd172;
	sample_rom[221][20] = 8'd156;
	sample_rom[221][21] = 8'd144;
	sample_rom[221][22] = 8'd141;
	sample_rom[221][23] = 8'd144;
	sample_rom[221][24] = 8'd150;
	sample_rom[221][25] = 8'd150;
	sample_rom[221][26] = 8'd144;
	sample_rom[221][27] = 8'd134;
	sample_rom[221][28] = 8'd116;
	sample_rom[221][29] = 8'd98;
	sample_rom[221][30] = 8'd83;
	sample_rom[221][31] = 8'd73;
	sample_rom[221][32] = 8'd73;
	sample_rom[221][33] = 8'd81;
	sample_rom[221][34] = 8'd94;
	sample_rom[221][35] = 8'd107;
	sample_rom[221][36] = 8'd119;
	sample_rom[221][37] = 8'd123;
	sample_rom[221][38] = 8'd117;
	sample_rom[221][39] = 8'd105;
	sample_rom[221][40] = 8'd90;
	sample_rom[221][41] = 8'd75;
	sample_rom[221][42] = 8'd63;
	sample_rom[221][43] = 8'd58;
	sample_rom[221][44] = 8'd60;
	sample_rom[221][45] = 8'd74;
	sample_rom[221][46] = 8'd87;
	sample_rom[221][47] = 8'd103;
	sample_rom[221][48] = 8'd115;
	sample_rom[221][49] = 8'd124;
	sample_rom[221][50] = 8'd126;
	sample_rom[221][51] = 8'd119;
	sample_rom[221][52] = 8'd114;
	sample_rom[221][53] = 8'd99;
	sample_rom[221][54] = 8'd95;
	sample_rom[221][55] = 8'd89;
	sample_rom[221][56] = 8'd91;
	sample_rom[221][57] = 8'd96;
	sample_rom[221][58] = 8'd103;
	sample_rom[221][59] = 8'd114;
	sample_rom[221][60] = 8'd124;
	sample_rom[221][61] = 8'd129;
	sample_rom[221][62] = 8'd134;
	sample_rom[221][63] = 8'd132;
	sample_rom[222][0] = 8'd131;
	sample_rom[222][1] = 8'd169;
	sample_rom[222][2] = 8'd202;
	sample_rom[222][3] = 8'd218;
	sample_rom[222][4] = 8'd218;
	sample_rom[222][5] = 8'd203;
	sample_rom[222][6] = 8'd182;
	sample_rom[222][7] = 8'd162;
	sample_rom[222][8] = 8'd153;
	sample_rom[222][9] = 8'd150;
	sample_rom[222][10] = 8'd158;
	sample_rom[222][11] = 8'd172;
	sample_rom[222][12] = 8'd187;
	sample_rom[222][13] = 8'd196;
	sample_rom[222][14] = 8'd197;
	sample_rom[222][15] = 8'd188;
	sample_rom[222][16] = 8'd171;
	sample_rom[222][17] = 8'd154;
	sample_rom[222][18] = 8'd139;
	sample_rom[222][19] = 8'd128;
	sample_rom[222][20] = 8'd124;
	sample_rom[222][21] = 8'd127;
	sample_rom[222][22] = 8'd127;
	sample_rom[222][23] = 8'd129;
	sample_rom[222][24] = 8'd121;
	sample_rom[222][25] = 8'd111;
	sample_rom[222][26] = 8'd97;
	sample_rom[222][27] = 8'd85;
	sample_rom[222][28] = 8'd78;
	sample_rom[222][29] = 8'd79;
	sample_rom[222][30] = 8'd89;
	sample_rom[222][31] = 8'd105;
	sample_rom[222][32] = 8'd124;
	sample_rom[222][33] = 8'd140;
	sample_rom[222][34] = 8'd151;
	sample_rom[222][35] = 8'd154;
	sample_rom[222][36] = 8'd150;
	sample_rom[222][37] = 8'd139;
	sample_rom[222][38] = 8'd131;
	sample_rom[222][39] = 8'd122;
	sample_rom[222][40] = 8'd118;
	sample_rom[222][41] = 8'd121;
	sample_rom[222][42] = 8'd124;
	sample_rom[222][43] = 8'd131;
	sample_rom[222][44] = 8'd134;
	sample_rom[222][45] = 8'd135;
	sample_rom[222][46] = 8'd131;
	sample_rom[222][47] = 8'd121;
	sample_rom[222][48] = 8'd110;
	sample_rom[222][49] = 8'd102;
	sample_rom[222][50] = 8'd97;
	sample_rom[222][51] = 8'd95;
	sample_rom[222][52] = 8'd96;
	sample_rom[222][53] = 8'd99;
	sample_rom[222][54] = 8'd103;
	sample_rom[222][55] = 8'd103;
	sample_rom[222][56] = 8'd102;
	sample_rom[222][57] = 8'd98;
	sample_rom[222][58] = 8'd93;
	sample_rom[222][59] = 8'd88;
	sample_rom[222][60] = 8'd87;
	sample_rom[222][61] = 8'd89;
	sample_rom[222][62] = 8'd99;
	sample_rom[222][63] = 8'd112;
	sample_rom[223][0] = 8'd131;
	sample_rom[223][1] = 8'd184;
	sample_rom[223][2] = 8'd219;
	sample_rom[223][3] = 8'd232;
	sample_rom[223][4] = 8'd221;
	sample_rom[223][5] = 8'd194;
	sample_rom[223][6] = 8'd165;
	sample_rom[223][7] = 8'd148;
	sample_rom[223][8] = 8'd149;
	sample_rom[223][9] = 8'd160;
	sample_rom[223][10] = 8'd181;
	sample_rom[223][11] = 8'd194;
	sample_rom[223][12] = 8'd198;
	sample_rom[223][13] = 8'd184;
	sample_rom[223][14] = 8'd162;
	sample_rom[223][15] = 8'd140;
	sample_rom[223][16] = 8'd118;
	sample_rom[223][17] = 8'd108;
	sample_rom[223][18] = 8'd105;
	sample_rom[223][19] = 8'd100;
	sample_rom[223][20] = 8'd97;
	sample_rom[223][21] = 8'd90;
	sample_rom[223][22] = 8'd79;
	sample_rom[223][23] = 8'd73;
	sample_rom[223][24] = 8'd72;
	sample_rom[223][25] = 8'd83;
	sample_rom[223][26] = 8'd103;
	sample_rom[223][27] = 8'd128;
	sample_rom[223][28] = 8'd149;
	sample_rom[223][29] = 8'd163;
	sample_rom[223][30] = 8'd165;
	sample_rom[223][31] = 8'd158;
	sample_rom[223][32] = 8'd144;
	sample_rom[223][33] = 8'd133;
	sample_rom[223][34] = 8'd128;
	sample_rom[223][35] = 8'd135;
	sample_rom[223][36] = 8'd145;
	sample_rom[223][37] = 8'd160;
	sample_rom[223][38] = 8'd174;
	sample_rom[223][39] = 8'd175;
	sample_rom[223][40] = 8'd172;
	sample_rom[223][41] = 8'd160;
	sample_rom[223][42] = 8'd145;
	sample_rom[223][43] = 8'd132;
	sample_rom[223][44] = 8'd124;
	sample_rom[223][45] = 8'd120;
	sample_rom[223][46] = 8'd120;
	sample_rom[223][47] = 8'd123;
	sample_rom[223][48] = 8'd125;
	sample_rom[223][49] = 8'd123;
	sample_rom[223][50] = 8'd125;
	sample_rom[223][51] = 8'd122;
	sample_rom[223][52] = 8'd125;
	sample_rom[223][53] = 8'd134;
	sample_rom[223][54] = 8'd143;
	sample_rom[223][55] = 8'd155;
	sample_rom[223][56] = 8'd159;
	sample_rom[223][57] = 8'd158;
	sample_rom[223][58] = 8'd149;
	sample_rom[223][59] = 8'd134;
	sample_rom[223][60] = 8'd119;
	sample_rom[223][61] = 8'd110;
	sample_rom[223][62] = 8'd109;
	sample_rom[223][63] = 8'd116;
	sample_rom[224][0] = 8'd130;
	sample_rom[224][1] = 8'd189;
	sample_rom[224][2] = 8'd225;
	sample_rom[224][3] = 8'd234;
	sample_rom[224][4] = 8'd220;
	sample_rom[224][5] = 8'd195;
	sample_rom[224][6] = 8'd173;
	sample_rom[224][7] = 8'd167;
	sample_rom[224][8] = 8'd177;
	sample_rom[224][9] = 8'd201;
	sample_rom[224][10] = 8'd215;
	sample_rom[224][11] = 8'd220;
	sample_rom[224][12] = 8'd209;
	sample_rom[224][13] = 8'd185;
	sample_rom[224][14] = 8'd164;
	sample_rom[224][15] = 8'd145;
	sample_rom[224][16] = 8'd134;
	sample_rom[224][17] = 8'd125;
	sample_rom[224][18] = 8'd112;
	sample_rom[224][19] = 8'd98;
	sample_rom[224][20] = 8'd83;
	sample_rom[224][21] = 8'd75;
	sample_rom[224][22] = 8'd76;
	sample_rom[224][23] = 8'd90;
	sample_rom[224][24] = 8'd110;
	sample_rom[224][25] = 8'd129;
	sample_rom[224][26] = 8'd140;
	sample_rom[224][27] = 8'd140;
	sample_rom[224][28] = 8'd129;
	sample_rom[224][29] = 8'd117;
	sample_rom[224][30] = 8'd113;
	sample_rom[224][31] = 8'd117;
	sample_rom[224][32] = 8'd126;
	sample_rom[224][33] = 8'd141;
	sample_rom[224][34] = 8'd151;
	sample_rom[224][35] = 8'd158;
	sample_rom[224][36] = 8'd155;
	sample_rom[224][37] = 8'd147;
	sample_rom[224][38] = 8'd142;
	sample_rom[224][39] = 8'd135;
	sample_rom[224][40] = 8'd129;
	sample_rom[224][41] = 8'd123;
	sample_rom[224][42] = 8'd118;
	sample_rom[224][43] = 8'd111;
	sample_rom[224][44] = 8'd109;
	sample_rom[224][45] = 8'd109;
	sample_rom[224][46] = 8'd121;
	sample_rom[224][47] = 8'd135;
	sample_rom[224][48] = 8'd151;
	sample_rom[224][49] = 8'd165;
	sample_rom[224][50] = 8'd172;
	sample_rom[224][51] = 8'd171;
	sample_rom[224][52] = 8'd167;
	sample_rom[224][53] = 8'd162;
	sample_rom[224][54] = 8'd160;
	sample_rom[224][55] = 8'd161;
	sample_rom[224][56] = 8'd170;
	sample_rom[224][57] = 8'd175;
	sample_rom[224][58] = 8'd182;
	sample_rom[224][59] = 8'd184;
	sample_rom[224][60] = 8'd177;
	sample_rom[224][61] = 8'd167;
	sample_rom[224][62] = 8'd156;
	sample_rom[224][63] = 8'd142;
	sample_rom[225][0] = 8'd131;
	sample_rom[225][1] = 8'd208;
	sample_rom[225][2] = 8'd250;
	sample_rom[225][3] = 8'd251;
	sample_rom[225][4] = 8'd221;
	sample_rom[225][5] = 8'd184;
	sample_rom[225][6] = 8'd169;
	sample_rom[225][7] = 8'd182;
	sample_rom[225][8] = 8'd210;
	sample_rom[225][9] = 8'd227;
	sample_rom[225][10] = 8'd227;
	sample_rom[225][11] = 8'd203;
	sample_rom[225][12] = 8'd171;
	sample_rom[225][13] = 8'd144;
	sample_rom[225][14] = 8'd130;
	sample_rom[225][15] = 8'd127;
	sample_rom[225][16] = 8'd117;
	sample_rom[225][17] = 8'd101;
	sample_rom[225][18] = 8'd83;
	sample_rom[225][19] = 8'd67;
	sample_rom[225][20] = 8'd71;
	sample_rom[225][21] = 8'd94;
	sample_rom[225][22] = 8'd126;
	sample_rom[225][23] = 8'd154;
	sample_rom[225][24] = 8'd164;
	sample_rom[225][25] = 8'd158;
	sample_rom[225][26] = 8'd142;
	sample_rom[225][27] = 8'd129;
	sample_rom[225][28] = 8'd128;
	sample_rom[225][29] = 8'd141;
	sample_rom[225][30] = 8'd152;
	sample_rom[225][31] = 8'd160;
	sample_rom[225][32] = 8'd157;
	sample_rom[225][33] = 8'd150;
	sample_rom[225][34] = 8'd136;
	sample_rom[225][35] = 8'd128;
	sample_rom[225][36] = 8'd121;
	sample_rom[225][37] = 8'd114;
	sample_rom[225][38] = 8'd108;
	sample_rom[225][39] = 8'd99;
	sample_rom[225][40] = 8'd97;
	sample_rom[225][41] = 8'd97;
	sample_rom[225][42] = 8'd111;
	sample_rom[225][43] = 8'd130;
	sample_rom[225][44] = 8'd152;
	sample_rom[225][45] = 8'd166;
	sample_rom[225][46] = 8'd173;
	sample_rom[225][47] = 8'd171;
	sample_rom[225][48] = 8'd167;
	sample_rom[225][49] = 8'd157;
	sample_rom[225][50] = 8'd158;
	sample_rom[225][51] = 8'd158;
	sample_rom[225][52] = 8'd166;
	sample_rom[225][53] = 8'd174;
	sample_rom[225][54] = 8'd177;
	sample_rom[225][55] = 8'd175;
	sample_rom[225][56] = 8'd169;
	sample_rom[225][57] = 8'd160;
	sample_rom[225][58] = 8'd146;
	sample_rom[225][59] = 8'd136;
	sample_rom[225][60] = 8'd124;
	sample_rom[225][61] = 8'd120;
	sample_rom[225][62] = 8'd121;
	sample_rom[225][63] = 8'd123;
	sample_rom[226][0] = 8'd129;
	sample_rom[226][1] = 8'd212;
	sample_rom[226][2] = 8'd249;
	sample_rom[226][3] = 8'd226;
	sample_rom[226][4] = 8'd176;
	sample_rom[226][5] = 8'd145;
	sample_rom[226][6] = 8'd148;
	sample_rom[226][7] = 8'd179;
	sample_rom[226][8] = 8'd204;
	sample_rom[226][9] = 8'd202;
	sample_rom[226][10] = 8'd177;
	sample_rom[226][11] = 8'd136;
	sample_rom[226][12] = 8'd117;
	sample_rom[226][13] = 8'd109;
	sample_rom[226][14] = 8'd105;
	sample_rom[226][15] = 8'd93;
	sample_rom[226][16] = 8'd67;
	sample_rom[226][17] = 8'd49;
	sample_rom[226][18] = 8'd52;
	sample_rom[226][19] = 8'd81;
	sample_rom[226][20] = 8'd115;
	sample_rom[226][21] = 8'd139;
	sample_rom[226][22] = 8'd139;
	sample_rom[226][23] = 8'd131;
	sample_rom[226][24] = 8'd121;
	sample_rom[226][25] = 8'd124;
	sample_rom[226][26] = 8'd140;
	sample_rom[226][27] = 8'd160;
	sample_rom[226][28] = 8'd164;
	sample_rom[226][29] = 8'd162;
	sample_rom[226][30] = 8'd152;
	sample_rom[226][31] = 8'd141;
	sample_rom[226][32] = 8'd134;
	sample_rom[226][33] = 8'd133;
	sample_rom[226][34] = 8'd123;
	sample_rom[226][35] = 8'd113;
	sample_rom[226][36] = 8'd102;
	sample_rom[226][37] = 8'd96;
	sample_rom[226][38] = 8'd100;
	sample_rom[226][39] = 8'd112;
	sample_rom[226][40] = 8'd128;
	sample_rom[226][41] = 8'd142;
	sample_rom[226][42] = 8'd142;
	sample_rom[226][43] = 8'd141;
	sample_rom[226][44] = 8'd135;
	sample_rom[226][45] = 8'd137;
	sample_rom[226][46] = 8'd140;
	sample_rom[226][47] = 8'd147;
	sample_rom[226][48] = 8'd151;
	sample_rom[226][49] = 8'd151;
	sample_rom[226][50] = 8'd148;
	sample_rom[226][51] = 8'd139;
	sample_rom[226][52] = 8'd133;
	sample_rom[226][53] = 8'd129;
	sample_rom[226][54] = 8'd120;
	sample_rom[226][55] = 8'd109;
	sample_rom[226][56] = 8'd100;
	sample_rom[226][57] = 8'd96;
	sample_rom[226][58] = 8'd94;
	sample_rom[226][59] = 8'd101;
	sample_rom[226][60] = 8'd111;
	sample_rom[226][61] = 8'd119;
	sample_rom[226][62] = 8'd128;
	sample_rom[226][63] = 8'd129;
	sample_rom[227][0] = 8'd130;
	sample_rom[227][1] = 8'd212;
	sample_rom[227][2] = 8'd237;
	sample_rom[227][3] = 8'd204;
	sample_rom[227][4] = 8'd163;
	sample_rom[227][5] = 8'd158;
	sample_rom[227][6] = 8'd188;
	sample_rom[227][7] = 8'd220;
	sample_rom[227][8] = 8'd212;
	sample_rom[227][9] = 8'd177;
	sample_rom[227][10] = 8'd139;
	sample_rom[227][11] = 8'd127;
	sample_rom[227][12] = 8'd125;
	sample_rom[227][13] = 8'd112;
	sample_rom[227][14] = 8'd84;
	sample_rom[227][15] = 8'd61;
	sample_rom[227][16] = 8'd65;
	sample_rom[227][17] = 8'd97;
	sample_rom[227][18] = 8'd126;
	sample_rom[227][19] = 8'd130;
	sample_rom[227][20] = 8'd114;
	sample_rom[227][21] = 8'd100;
	sample_rom[227][22] = 8'd105;
	sample_rom[227][23] = 8'd127;
	sample_rom[227][24] = 8'd145;
	sample_rom[227][25] = 8'd144;
	sample_rom[227][26] = 8'd131;
	sample_rom[227][27] = 8'd119;
	sample_rom[227][28] = 8'd115;
	sample_rom[227][29] = 8'd120;
	sample_rom[227][30] = 8'd117;
	sample_rom[227][31] = 8'd104;
	sample_rom[227][32] = 8'd98;
	sample_rom[227][33] = 8'd103;
	sample_rom[227][34] = 8'd122;
	sample_rom[227][35] = 8'd143;
	sample_rom[227][36] = 8'd157;
	sample_rom[227][37] = 8'd154;
	sample_rom[227][38] = 8'd149;
	sample_rom[227][39] = 8'd148;
	sample_rom[227][40] = 8'd157;
	sample_rom[227][41] = 8'd168;
	sample_rom[227][42] = 8'd171;
	sample_rom[227][43] = 8'd167;
	sample_rom[227][44] = 8'd153;
	sample_rom[227][45] = 8'd143;
	sample_rom[227][46] = 8'd135;
	sample_rom[227][47] = 8'd129;
	sample_rom[227][48] = 8'd119;
	sample_rom[227][49] = 8'd102;
	sample_rom[227][50] = 8'd93;
	sample_rom[227][51] = 8'd94;
	sample_rom[227][52] = 8'd103;
	sample_rom[227][53] = 8'd113;
	sample_rom[227][54] = 8'd115;
	sample_rom[227][55] = 8'd106;
	sample_rom[227][56] = 8'd99;
	sample_rom[227][57] = 8'd102;
	sample_rom[227][58] = 8'd111;
	sample_rom[227][59] = 8'd126;
	sample_rom[227][60] = 8'd131;
	sample_rom[227][61] = 8'd132;
	sample_rom[227][62] = 8'd128;
	sample_rom[227][63] = 8'd126;
	sample_rom[228][0] = 8'd130;
	sample_rom[228][1] = 8'd226;
	sample_rom[228][2] = 8'd245;
	sample_rom[228][3] = 8'd198;
	sample_rom[228][4] = 8'd156;
	sample_rom[228][5] = 8'd167;
	sample_rom[228][6] = 8'd207;
	sample_rom[228][7] = 8'd223;
	sample_rom[228][8] = 8'd186;
	sample_rom[228][9] = 8'd143;
	sample_rom[228][10] = 8'd118;
	sample_rom[228][11] = 8'd119;
	sample_rom[228][12] = 8'd106;
	sample_rom[228][13] = 8'd74;
	sample_rom[228][14] = 8'd52;
	sample_rom[228][15] = 8'd70;
	sample_rom[228][16] = 8'd112;
	sample_rom[228][17] = 8'd139;
	sample_rom[228][18] = 8'd137;
	sample_rom[228][19] = 8'd118;
	sample_rom[228][20] = 8'd116;
	sample_rom[228][21] = 8'd134;
	sample_rom[228][22] = 8'd156;
	sample_rom[228][23] = 8'd152;
	sample_rom[228][24] = 8'd132;
	sample_rom[228][25] = 8'd117;
	sample_rom[228][26] = 8'd117;
	sample_rom[228][27] = 8'd117;
	sample_rom[228][28] = 8'd105;
	sample_rom[228][29] = 8'd90;
	sample_rom[228][30] = 8'd84;
	sample_rom[228][31] = 8'd97;
	sample_rom[228][32] = 8'd123;
	sample_rom[228][33] = 8'd145;
	sample_rom[228][34] = 8'd148;
	sample_rom[228][35] = 8'd146;
	sample_rom[228][36] = 8'd147;
	sample_rom[228][37] = 8'd157;
	sample_rom[228][38] = 8'd165;
	sample_rom[228][39] = 8'd165;
	sample_rom[228][40] = 8'd157;
	sample_rom[228][41] = 8'd148;
	sample_rom[228][42] = 8'd144;
	sample_rom[228][43] = 8'd144;
	sample_rom[228][44] = 8'd127;
	sample_rom[228][45] = 8'd113;
	sample_rom[228][46] = 8'd103;
	sample_rom[228][47] = 8'd104;
	sample_rom[228][48] = 8'd119;
	sample_rom[228][49] = 8'd128;
	sample_rom[228][50] = 8'd128;
	sample_rom[228][51] = 8'd120;
	sample_rom[228][52] = 8'd115;
	sample_rom[228][53] = 8'd120;
	sample_rom[228][54] = 8'd124;
	sample_rom[228][55] = 8'd124;
	sample_rom[228][56] = 8'd121;
	sample_rom[228][57] = 8'd118;
	sample_rom[228][58] = 8'd118;
	sample_rom[228][59] = 8'd121;
	sample_rom[228][60] = 8'd118;
	sample_rom[228][61] = 8'd114;
	sample_rom[228][62] = 8'd111;
	sample_rom[228][63] = 8'd116;
	sample_rom[229][0] = 8'd128;
	sample_rom[229][1] = 8'd220;
	sample_rom[229][2] = 8'd220;
	sample_rom[229][3] = 8'd167;
	sample_rom[229][4] = 8'd156;
	sample_rom[229][5] = 8'd188;
	sample_rom[229][6] = 8'd205;
	sample_rom[229][7] = 8'd169;
	sample_rom[229][8] = 8'd131;
	sample_rom[229][9] = 8'd118;
	sample_rom[229][10] = 8'd109;
	sample_rom[229][11] = 8'd84;
	sample_rom[229][12] = 8'd66;
	sample_rom[229][13] = 8'd99;
	sample_rom[229][14] = 8'd141;
	sample_rom[229][15] = 8'd153;
	sample_rom[229][16] = 8'd128;
	sample_rom[229][17] = 8'd119;
	sample_rom[229][18] = 8'd138;
	sample_rom[229][19] = 8'd155;
	sample_rom[229][20] = 8'd147;
	sample_rom[229][21] = 8'd128;
	sample_rom[229][22] = 8'd117;
	sample_rom[229][23] = 8'd116;
	sample_rom[229][24] = 8'd108;
	sample_rom[229][25] = 8'd103;
	sample_rom[229][26] = 8'd113;
	sample_rom[229][27] = 8'd140;
	sample_rom[229][28] = 8'd159;
	sample_rom[229][29] = 8'd151;
	sample_rom[229][30] = 8'd141;
	sample_rom[229][31] = 8'd143;
	sample_rom[229][32] = 8'd156;
	sample_rom[229][33] = 8'd159;
	sample_rom[229][34] = 8'd147;
	sample_rom[229][35] = 8'd133;
	sample_rom[229][36] = 8'd128;
	sample_rom[229][37] = 8'd124;
	sample_rom[229][38] = 8'd114;
	sample_rom[229][39] = 8'd106;
	sample_rom[229][40] = 8'd114;
	sample_rom[229][41] = 8'd122;
	sample_rom[229][42] = 8'd123;
	sample_rom[229][43] = 8'd109;
	sample_rom[229][44] = 8'd104;
	sample_rom[229][45] = 8'd111;
	sample_rom[229][46] = 8'd119;
	sample_rom[229][47] = 8'd116;
	sample_rom[229][48] = 8'd115;
	sample_rom[229][49] = 8'd115;
	sample_rom[229][50] = 8'd119;
	sample_rom[229][51] = 8'd121;
	sample_rom[229][52] = 8'd125;
	sample_rom[229][53] = 8'd129;
	sample_rom[229][54] = 8'd139;
	sample_rom[229][55] = 8'd143;
	sample_rom[229][56] = 8'd136;
	sample_rom[229][57] = 8'd135;
	sample_rom[229][58] = 8'd134;
	sample_rom[229][59] = 8'd136;
	sample_rom[229][60] = 8'd135;
	sample_rom[229][61] = 8'd130;
	sample_rom[229][62] = 8'd127;
	sample_rom[229][63] = 8'd128;
	sample_rom[230][0] = 8'd128;
	sample_rom[230][1] = 8'd221;
	sample_rom[230][2] = 8'd221;
	sample_rom[230][3] = 8'd171;
	sample_rom[230][4] = 8'd170;
	sample_rom[230][5] = 8'd202;
	sample_rom[230][6] = 8'd198;
	sample_rom[230][7] = 8'd147;
	sample_rom[230][8] = 8'd115;
	sample_rom[230][9] = 8'd104;
	sample_rom[230][10] = 8'd86;
	sample_rom[230][11] = 8'd72;
	sample_rom[230][12] = 8'd99;
	sample_rom[230][13] = 8'd142;
	sample_rom[230][14] = 8'd146;
	sample_rom[230][15] = 8'd125;
	sample_rom[230][16] = 8'd124;
	sample_rom[230][17] = 8'd156;
	sample_rom[230][18] = 8'd159;
	sample_rom[230][19] = 8'd134;
	sample_rom[230][20] = 8'd117;
	sample_rom[230][21] = 8'd119;
	sample_rom[230][22] = 8'd113;
	sample_rom[230][23] = 8'd107;
	sample_rom[230][24] = 8'd126;
	sample_rom[230][25] = 8'd159;
	sample_rom[230][26] = 8'd164;
	sample_rom[230][27] = 8'd147;
	sample_rom[230][28] = 8'd140;
	sample_rom[230][29] = 8'd160;
	sample_rom[230][30] = 8'd162;
	sample_rom[230][31] = 8'd143;
	sample_rom[230][32] = 8'd123;
	sample_rom[230][33] = 8'd119;
	sample_rom[230][34] = 8'd112;
	sample_rom[230][35] = 8'd103;
	sample_rom[230][36] = 8'd105;
	sample_rom[230][37] = 8'd120;
	sample_rom[230][38] = 8'd123;
	sample_rom[230][39] = 8'd110;
	sample_rom[230][40] = 8'd103;
	sample_rom[230][41] = 8'd119;
	sample_rom[230][42] = 8'd131;
	sample_rom[230][43] = 8'd126;
	sample_rom[230][44] = 8'd120;
	sample_rom[230][45] = 8'd123;
	sample_rom[230][46] = 8'd127;
	sample_rom[230][47] = 8'd130;
	sample_rom[230][48] = 8'd130;
	sample_rom[230][49] = 8'd137;
	sample_rom[230][50] = 8'd141;
	sample_rom[230][51] = 8'd130;
	sample_rom[230][52] = 8'd119;
	sample_rom[230][53] = 8'd120;
	sample_rom[230][54] = 8'd123;
	sample_rom[230][55] = 8'd120;
	sample_rom[230][56] = 8'd112;
	sample_rom[230][57] = 8'd115;
	sample_rom[230][58] = 8'd115;
	sample_rom[230][59] = 8'd119;
	sample_rom[230][60] = 8'd122;
	sample_rom[230][61] = 8'd124;
	sample_rom[230][62] = 8'd127;
	sample_rom[230][63] = 8'd130;
	sample_rom[231][0] = 8'd128;
	sample_rom[231][1] = 8'd208;
	sample_rom[231][2] = 8'd216;
	sample_rom[231][3] = 8'd185;
	sample_rom[231][4] = 8'd179;
	sample_rom[231][5] = 8'd195;
	sample_rom[231][6] = 8'd183;
	sample_rom[231][7] = 8'd131;
	sample_rom[231][8] = 8'd86;
	sample_rom[231][9] = 8'd77;
	sample_rom[231][10] = 8'd93;
	sample_rom[231][11] = 8'd114;
	sample_rom[231][12] = 8'd126;
	sample_rom[231][13] = 8'd137;
	sample_rom[231][14] = 8'd143;
	sample_rom[231][15] = 8'd144;
	sample_rom[231][16] = 8'd149;
	sample_rom[231][17] = 8'd147;
	sample_rom[231][18] = 8'd128;
	sample_rom[231][19] = 8'd102;
	sample_rom[231][20] = 8'd101;
	sample_rom[231][21] = 8'd120;
	sample_rom[231][22] = 8'd141;
	sample_rom[231][23] = 8'd152;
	sample_rom[231][24] = 8'd153;
	sample_rom[231][25] = 8'd161;
	sample_rom[231][26] = 8'd163;
	sample_rom[231][27] = 8'd161;
	sample_rom[231][28] = 8'd153;
	sample_rom[231][29] = 8'd137;
	sample_rom[231][30] = 8'd114;
	sample_rom[231][31] = 8'd105;
	sample_rom[231][32] = 8'd108;
	sample_rom[231][33] = 8'd117;
	sample_rom[231][34] = 8'd117;
	sample_rom[231][35] = 8'd115;
	sample_rom[231][36] = 8'd110;
	sample_rom[231][37] = 8'd121;
	sample_rom[231][38] = 8'd127;
	sample_rom[231][39] = 8'd124;
	sample_rom[231][40] = 8'd118;
	sample_rom[231][41] = 8'd114;
	sample_rom[231][42] = 8'd119;
	sample_rom[231][43] = 8'd128;
	sample_rom[231][44] = 8'd137;
	sample_rom[231][45] = 8'd137;
	sample_rom[231][46] = 8'd130;
	sample_rom[231][47] = 8'd126;
	sample_rom[231][48] = 8'd128;
	sample_rom[231][49] = 8'd133;
	sample_rom[231][50] = 8'd124;
	sample_rom[231][51] = 8'd113;
	sample_rom[231][52] = 8'd112;
	sample_rom[231][53] = 8'd117;
	sample_rom[231][54] = 8'd124;
	sample_rom[231][55] = 8'd127;
	sample_rom[231][56] = 8'd123;
	sample_rom[231][57] = 8'd119;
	sample_rom[231][58] = 8'd116;
	sample_rom[231][59] = 8'd119;
	sample_rom[231][60] = 8'd119;
	sample_rom[231][61] = 8'd117;
	sample_rom[231][62] = 8'd115;
	sample_rom[231][63] = 8'd117;
	sample_rom[232][0] = 8'd128;
	sample_rom[232][1] = 8'd212;
	sample_rom[232][2] = 8'd218;
	sample_rom[232][3] = 8'd186;
	sample_rom[232][4] = 8'd179;
	sample_rom[232][5] = 8'd190;
	sample_rom[232][6] = 8'd157;
	sample_rom[232][7] = 8'd89;
	sample_rom[232][8] = 8'd54;
	sample_rom[232][9] = 8'd76;
	sample_rom[232][10] = 8'd114;
	sample_rom[232][11] = 8'd124;
	sample_rom[232][12] = 8'd120;
	sample_rom[232][13] = 8'd131;
	sample_rom[232][14] = 8'd148;
	sample_rom[232][15] = 8'd146;
	sample_rom[232][16] = 8'd124;
	sample_rom[232][17] = 8'd103;
	sample_rom[232][18] = 8'd99;
	sample_rom[232][19] = 8'd113;
	sample_rom[232][20] = 8'd137;
	sample_rom[232][21] = 8'd151;
	sample_rom[232][22] = 8'd153;
	sample_rom[232][23] = 8'd154;
	sample_rom[232][24] = 8'd160;
	sample_rom[232][25] = 8'd159;
	sample_rom[232][26] = 8'd141;
	sample_rom[232][27] = 8'd110;
	sample_rom[232][28] = 8'd99;
	sample_rom[232][29] = 8'd109;
	sample_rom[232][30] = 8'd116;
	sample_rom[232][31] = 8'd110;
	sample_rom[232][32] = 8'd108;
	sample_rom[232][33] = 8'd119;
	sample_rom[232][34] = 8'd132;
	sample_rom[232][35] = 8'd135;
	sample_rom[232][36] = 8'd129;
	sample_rom[232][37] = 8'd126;
	sample_rom[232][38] = 8'd130;
	sample_rom[232][39] = 8'd138;
	sample_rom[232][40] = 8'd145;
	sample_rom[232][41] = 8'd143;
	sample_rom[232][42] = 8'd138;
	sample_rom[232][43] = 8'd136;
	sample_rom[232][44] = 8'd139;
	sample_rom[232][45] = 8'd136;
	sample_rom[232][46] = 8'd123;
	sample_rom[232][47] = 8'd112;
	sample_rom[232][48] = 8'd112;
	sample_rom[232][49] = 8'd119;
	sample_rom[232][50] = 8'd121;
	sample_rom[232][51] = 8'd116;
	sample_rom[232][52] = 8'd119;
	sample_rom[232][53] = 8'd126;
	sample_rom[232][54] = 8'd132;
	sample_rom[232][55] = 8'd129;
	sample_rom[232][56] = 8'd129;
	sample_rom[232][57] = 8'd134;
	sample_rom[232][58] = 8'd140;
	sample_rom[232][59] = 8'd143;
	sample_rom[232][60] = 8'd142;
	sample_rom[232][61] = 8'd142;
	sample_rom[232][62] = 8'd140;
	sample_rom[232][63] = 8'd136;
	sample_rom[233][0] = 8'd128;
	sample_rom[233][1] = 8'd212;
	sample_rom[233][2] = 8'd228;
	sample_rom[233][3] = 8'd209;
	sample_rom[233][4] = 8'd193;
	sample_rom[233][5] = 8'd167;
	sample_rom[233][6] = 8'd109;
	sample_rom[233][7] = 8'd59;
	sample_rom[233][8] = 8'd70;
	sample_rom[233][9] = 8'd118;
	sample_rom[233][10] = 8'd138;
	sample_rom[233][11] = 8'd133;
	sample_rom[233][12] = 8'd145;
	sample_rom[233][13] = 8'd159;
	sample_rom[233][14] = 8'd138;
	sample_rom[233][15] = 8'd99;
	sample_rom[233][16] = 8'd98;
	sample_rom[233][17] = 8'd137;
	sample_rom[233][18] = 8'd159;
	sample_rom[233][19] = 8'd154;
	sample_rom[233][20] = 8'd156;
	sample_rom[233][21] = 8'd168;
	sample_rom[233][22] = 8'd158;
	sample_rom[233][23] = 8'd118;
	sample_rom[233][24] = 8'd90;
	sample_rom[233][25] = 8'd98;
	sample_rom[233][26] = 8'd109;
	sample_rom[233][27] = 8'd102;
	sample_rom[233][28] = 8'd101;
	sample_rom[233][29] = 8'd122;
	sample_rom[233][30] = 8'd136;
	sample_rom[233][31] = 8'd125;
	sample_rom[233][32] = 8'd113;
	sample_rom[233][33] = 8'd123;
	sample_rom[233][34] = 8'd138;
	sample_rom[233][35] = 8'd135;
	sample_rom[233][36] = 8'd130;
	sample_rom[233][37] = 8'd135;
	sample_rom[233][38] = 8'd137;
	sample_rom[233][39] = 8'd128;
	sample_rom[233][40] = 8'd114;
	sample_rom[233][41] = 8'd110;
	sample_rom[233][42] = 8'd117;
	sample_rom[233][43] = 8'd120;
	sample_rom[233][44] = 8'd121;
	sample_rom[233][45] = 8'd124;
	sample_rom[233][46] = 8'd131;
	sample_rom[233][47] = 8'd135;
	sample_rom[233][48] = 8'd134;
	sample_rom[233][49] = 8'd134;
	sample_rom[233][50] = 8'd140;
	sample_rom[233][51] = 8'd146;
	sample_rom[233][52] = 8'd150;
	sample_rom[233][53] = 8'd149;
	sample_rom[233][54] = 8'd146;
	sample_rom[233][55] = 8'd138;
	sample_rom[233][56] = 8'd133;
	sample_rom[233][57] = 8'd127;
	sample_rom[233][58] = 8'd121;
	sample_rom[233][59] = 8'd119;
	sample_rom[233][60] = 8'd124;
	sample_rom[233][61] = 8'd128;
	sample_rom[233][62] = 8'd128;
	sample_rom[233][63] = 8'd126;
	sample_rom[234][0] = 8'd128;
	sample_rom[234][1] = 8'd208;
	sample_rom[234][2] = 8'd238;
	sample_rom[234][3] = 8'd223;
	sample_rom[234][4] = 8'd188;
	sample_rom[234][5] = 8'd135;
	sample_rom[234][6] = 8'd84;
	sample_rom[234][7] = 8'd62;
	sample_rom[234][8] = 8'd86;
	sample_rom[234][9] = 8'd125;
	sample_rom[234][10] = 8'd144;
	sample_rom[234][11] = 8'd143;
	sample_rom[234][12] = 8'd140;
	sample_rom[234][13] = 8'd125;
	sample_rom[234][14] = 8'd103;
	sample_rom[234][15] = 8'd103;
	sample_rom[234][16] = 8'd128;
	sample_rom[234][17] = 8'd162;
	sample_rom[234][18] = 8'd172;
	sample_rom[234][19] = 8'd166;
	sample_rom[234][20] = 8'd160;
	sample_rom[234][21] = 8'd145;
	sample_rom[234][22] = 8'd115;
	sample_rom[234][23] = 8'd95;
	sample_rom[234][24] = 8'd98;
	sample_rom[234][25] = 8'd110;
	sample_rom[234][26] = 8'd112;
	sample_rom[234][27] = 8'd112;
	sample_rom[234][28] = 8'd124;
	sample_rom[234][29] = 8'd129;
	sample_rom[234][30] = 8'd124;
	sample_rom[234][31] = 8'd120;
	sample_rom[234][32] = 8'd133;
	sample_rom[234][33] = 8'd145;
	sample_rom[234][34] = 8'd140;
	sample_rom[234][35] = 8'd130;
	sample_rom[234][36] = 8'd132;
	sample_rom[234][37] = 8'd130;
	sample_rom[234][38] = 8'd118;
	sample_rom[234][39] = 8'd107;
	sample_rom[234][40] = 8'd114;
	sample_rom[234][41] = 8'd124;
	sample_rom[234][42] = 8'd120;
	sample_rom[234][43] = 8'd117;
	sample_rom[234][44] = 8'd125;
	sample_rom[234][45] = 8'd136;
	sample_rom[234][46] = 8'd133;
	sample_rom[234][47] = 8'd134;
	sample_rom[234][48] = 8'd142;
	sample_rom[234][49] = 8'd151;
	sample_rom[234][50] = 8'd140;
	sample_rom[234][51] = 8'd130;
	sample_rom[234][52] = 8'd130;
	sample_rom[234][53] = 8'd134;
	sample_rom[234][54] = 8'd129;
	sample_rom[234][55] = 8'd121;
	sample_rom[234][56] = 8'd129;
	sample_rom[234][57] = 8'd137;
	sample_rom[234][58] = 8'd131;
	sample_rom[234][59] = 8'd125;
	sample_rom[234][60] = 8'd135;
	sample_rom[234][61] = 8'd140;
	sample_rom[234][62] = 8'd133;
	sample_rom[234][63] = 8'd125;
	sample_rom[235][0] = 8'd128;
	sample_rom[235][1] = 8'd209;
	sample_rom[235][2] = 8'd238;
	sample_rom[235][3] = 8'd209;
	sample_rom[235][4] = 8'd142;
	sample_rom[235][5] = 8'd87;
	sample_rom[235][6] = 8'd74;
	sample_rom[235][7] = 8'd99;
	sample_rom[235][8] = 8'd136;
	sample_rom[235][9] = 8'd157;
	sample_rom[235][10] = 8'd146;
	sample_rom[235][11] = 8'd123;
	sample_rom[235][12] = 8'd110;
	sample_rom[235][13] = 8'd121;
	sample_rom[235][14] = 8'd145;
	sample_rom[235][15] = 8'd170;
	sample_rom[235][16] = 8'd172;
	sample_rom[235][17] = 8'd150;
	sample_rom[235][18] = 8'd122;
	sample_rom[235][19] = 8'd105;
	sample_rom[235][20] = 8'd101;
	sample_rom[235][21] = 8'd108;
	sample_rom[235][22] = 8'd115;
	sample_rom[235][23] = 8'd119;
	sample_rom[235][24] = 8'd120;
	sample_rom[235][25] = 8'd123;
	sample_rom[235][26] = 8'd132;
	sample_rom[235][27] = 8'd141;
	sample_rom[235][28] = 8'd141;
	sample_rom[235][29] = 8'd134;
	sample_rom[235][30] = 8'd124;
	sample_rom[235][31] = 8'd113;
	sample_rom[235][32] = 8'd111;
	sample_rom[235][33] = 8'd114;
	sample_rom[235][34] = 8'd117;
	sample_rom[235][35] = 8'd120;
	sample_rom[235][36] = 8'd126;
	sample_rom[235][37] = 8'd128;
	sample_rom[235][38] = 8'd134;
	sample_rom[235][39] = 8'd139;
	sample_rom[235][40] = 8'd144;
	sample_rom[235][41] = 8'd143;
	sample_rom[235][42] = 8'd139;
	sample_rom[235][43] = 8'd129;
	sample_rom[235][44] = 8'd125;
	sample_rom[235][45] = 8'd122;
	sample_rom[235][46] = 8'd128;
	sample_rom[235][47] = 8'd128;
	sample_rom[235][48] = 8'd128;
	sample_rom[235][49] = 8'd127;
	sample_rom[235][50] = 8'd129;
	sample_rom[235][51] = 8'd133;
	sample_rom[235][52] = 8'd137;
	sample_rom[235][53] = 8'd139;
	sample_rom[235][54] = 8'd133;
	sample_rom[235][55] = 8'd124;
	sample_rom[235][56] = 8'd120;
	sample_rom[235][57] = 8'd120;
	sample_rom[235][58] = 8'd127;
	sample_rom[235][59] = 8'd132;
	sample_rom[235][60] = 8'd131;
	sample_rom[235][61] = 8'd127;
	sample_rom[235][62] = 8'd123;
	sample_rom[235][63] = 8'd123;
	sample_rom[236][0] = 8'd128;
	sample_rom[236][1] = 8'd222;
	sample_rom[236][2] = 8'd245;
	sample_rom[236][3] = 8'd196;
	sample_rom[236][4] = 8'd114;
	sample_rom[236][5] = 8'd67;
	sample_rom[236][6] = 8'd81;
	sample_rom[236][7] = 8'd125;
	sample_rom[236][8] = 8'd154;
	sample_rom[236][9] = 8'd147;
	sample_rom[236][10] = 8'd116;
	sample_rom[236][11] = 8'd100;
	sample_rom[236][12] = 8'd121;
	sample_rom[236][13] = 8'd155;
	sample_rom[236][14] = 8'd175;
	sample_rom[236][15] = 8'd166;
	sample_rom[236][16] = 8'd136;
	sample_rom[236][17] = 8'd108;
	sample_rom[236][18] = 8'd98;
	sample_rom[236][19] = 8'd105;
	sample_rom[236][20] = 8'd113;
	sample_rom[236][21] = 8'd120;
	sample_rom[236][22] = 8'd122;
	sample_rom[236][23] = 8'd124;
	sample_rom[236][24] = 8'd133;
	sample_rom[236][25] = 8'd144;
	sample_rom[236][26] = 8'd142;
	sample_rom[236][27] = 8'd132;
	sample_rom[236][28] = 8'd121;
	sample_rom[236][29] = 8'd115;
	sample_rom[236][30] = 8'd115;
	sample_rom[236][31] = 8'd120;
	sample_rom[236][32] = 8'd121;
	sample_rom[236][33] = 8'd125;
	sample_rom[236][34] = 8'd127;
	sample_rom[236][35] = 8'd135;
	sample_rom[236][36] = 8'd142;
	sample_rom[236][37] = 8'd149;
	sample_rom[236][38] = 8'd142;
	sample_rom[236][39] = 8'd132;
	sample_rom[236][40] = 8'd127;
	sample_rom[236][41] = 8'd126;
	sample_rom[236][42] = 8'd130;
	sample_rom[236][43] = 8'd131;
	sample_rom[236][44] = 8'd130;
	sample_rom[236][45] = 8'd131;
	sample_rom[236][46] = 8'd131;
	sample_rom[236][47] = 8'd133;
	sample_rom[236][48] = 8'd137;
	sample_rom[236][49] = 8'd134;
	sample_rom[236][50] = 8'd126;
	sample_rom[236][51] = 8'd120;
	sample_rom[236][52] = 8'd118;
	sample_rom[236][53] = 8'd123;
	sample_rom[236][54] = 8'd127;
	sample_rom[236][55] = 8'd126;
	sample_rom[236][56] = 8'd123;
	sample_rom[236][57] = 8'd123;
	sample_rom[236][58] = 8'd123;
	sample_rom[236][59] = 8'd127;
	sample_rom[236][60] = 8'd128;
	sample_rom[236][61] = 8'd125;
	sample_rom[236][62] = 8'd119;
	sample_rom[236][63] = 8'd122;
	sample_rom[237][0] = 8'd128;
	sample_rom[237][1] = 8'd239;
	sample_rom[237][2] = 8'd252;
	sample_rom[237][3] = 8'd170;
	sample_rom[237][4] = 8'd85;
	sample_rom[237][5] = 8'd63;
	sample_rom[237][6] = 8'd109;
	sample_rom[237][7] = 8'd156;
	sample_rom[237][8] = 8'd156;
	sample_rom[237][9] = 8'd122;
	sample_rom[237][10] = 8'd105;
	sample_rom[237][11] = 8'd129;
	sample_rom[237][12] = 8'd169;
	sample_rom[237][13] = 8'd183;
	sample_rom[237][14] = 8'd154;
	sample_rom[237][15] = 8'd110;
	sample_rom[237][16] = 8'd90;
	sample_rom[237][17] = 8'd97;
	sample_rom[237][18] = 8'd115;
	sample_rom[237][19] = 8'd122;
	sample_rom[237][20] = 8'd122;
	sample_rom[237][21] = 8'd125;
	sample_rom[237][22] = 8'd135;
	sample_rom[237][23] = 8'd142;
	sample_rom[237][24] = 8'd135;
	sample_rom[237][25] = 8'd120;
	sample_rom[237][26] = 8'd110;
	sample_rom[237][27] = 8'd108;
	sample_rom[237][28] = 8'd119;
	sample_rom[237][29] = 8'd125;
	sample_rom[237][30] = 8'd125;
	sample_rom[237][31] = 8'd130;
	sample_rom[237][32] = 8'd136;
	sample_rom[237][33] = 8'd146;
	sample_rom[237][34] = 8'd151;
	sample_rom[237][35] = 8'd139;
	sample_rom[237][36] = 8'd130;
	sample_rom[237][37] = 8'd120;
	sample_rom[237][38] = 8'd126;
	sample_rom[237][39] = 8'd133;
	sample_rom[237][40] = 8'd135;
	sample_rom[237][41] = 8'd134;
	sample_rom[237][42] = 8'd133;
	sample_rom[237][43] = 8'd136;
	sample_rom[237][44] = 8'd138;
	sample_rom[237][45] = 8'd133;
	sample_rom[237][46] = 8'd126;
	sample_rom[237][47] = 8'd122;
	sample_rom[237][48] = 8'd122;
	sample_rom[237][49] = 8'd127;
	sample_rom[237][50] = 8'd126;
	sample_rom[237][51] = 8'd123;
	sample_rom[237][52] = 8'd124;
	sample_rom[237][53] = 8'd125;
	sample_rom[237][54] = 8'd131;
	sample_rom[237][55] = 8'd133;
	sample_rom[237][56] = 8'd127;
	sample_rom[237][57] = 8'd123;
	sample_rom[237][58] = 8'd123;
	sample_rom[237][59] = 8'd124;
	sample_rom[237][60] = 8'd128;
	sample_rom[237][61] = 8'd128;
	sample_rom[237][62] = 8'd124;
	sample_rom[237][63] = 8'd127;
	sample_rom[238][0] = 8'd128;
	sample_rom[238][1] = 8'd207;
	sample_rom[238][2] = 8'd203;
	sample_rom[238][3] = 8'd132;
	sample_rom[238][4] = 8'd82;
	sample_rom[238][5] = 8'd97;
	sample_rom[238][6] = 8'd138;
	sample_rom[238][7] = 8'd146;
	sample_rom[238][8] = 8'd120;
	sample_rom[238][9] = 8'd110;
	sample_rom[238][10] = 8'd135;
	sample_rom[238][11] = 8'd162;
	sample_rom[238][12] = 8'd161;
	sample_rom[238][13] = 8'd133;
	sample_rom[238][14] = 8'd108;
	sample_rom[238][15] = 8'd106;
	sample_rom[238][16] = 8'd116;
	sample_rom[238][17] = 8'd122;
	sample_rom[238][18] = 8'd124;
	sample_rom[238][19] = 8'd130;
	sample_rom[238][20] = 8'd137;
	sample_rom[238][21] = 8'd139;
	sample_rom[238][22] = 8'd129;
	sample_rom[238][23] = 8'd119;
	sample_rom[238][24] = 8'd117;
	sample_rom[238][25] = 8'd121;
	sample_rom[238][26] = 8'd125;
	sample_rom[238][27] = 8'd128;
	sample_rom[238][28] = 8'd133;
	sample_rom[238][29] = 8'd138;
	sample_rom[238][30] = 8'd144;
	sample_rom[238][31] = 8'd136;
	sample_rom[238][32] = 8'd129;
	sample_rom[238][33] = 8'd126;
	sample_rom[238][34] = 8'd126;
	sample_rom[238][35] = 8'd128;
	sample_rom[238][36] = 8'd128;
	sample_rom[238][37] = 8'd128;
	sample_rom[238][38] = 8'd128;
	sample_rom[238][39] = 8'd133;
	sample_rom[238][40] = 8'd130;
	sample_rom[238][41] = 8'd127;
	sample_rom[238][42] = 8'd124;
	sample_rom[238][43] = 8'd124;
	sample_rom[238][44] = 8'd127;
	sample_rom[238][45] = 8'd124;
	sample_rom[238][46] = 8'd120;
	sample_rom[238][47] = 8'd123;
	sample_rom[238][48] = 8'd126;
	sample_rom[238][49] = 8'd129;
	sample_rom[238][50] = 8'd127;
	sample_rom[238][51] = 8'd127;
	sample_rom[238][52] = 8'd129;
	sample_rom[238][53] = 8'd134;
	sample_rom[238][54] = 8'd132;
	sample_rom[238][55] = 8'd131;
	sample_rom[238][56] = 8'd126;
	sample_rom[238][57] = 8'd128;
	sample_rom[238][58] = 8'd130;
	sample_rom[238][59] = 8'd132;
	sample_rom[238][60] = 8'd128;
	sample_rom[238][61] = 8'd131;
	sample_rom[238][62] = 8'd132;
	sample_rom[238][63] = 8'd134;
	sample_rom[239][0] = 8'd128;
	sample_rom[239][1] = 8'd207;
	sample_rom[239][2] = 8'd203;
	sample_rom[239][3] = 8'd132;
	sample_rom[239][4] = 8'd82;
	sample_rom[239][5] = 8'd97;
	sample_rom[239][6] = 8'd138;
	sample_rom[239][7] = 8'd146;
	sample_rom[239][8] = 8'd120;
	sample_rom[239][9] = 8'd110;
	sample_rom[239][10] = 8'd135;
	sample_rom[239][11] = 8'd162;
	sample_rom[239][12] = 8'd161;
	sample_rom[239][13] = 8'd133;
	sample_rom[239][14] = 8'd108;
	sample_rom[239][15] = 8'd106;
	sample_rom[239][16] = 8'd116;
	sample_rom[239][17] = 8'd122;
	sample_rom[239][18] = 8'd124;
	sample_rom[239][19] = 8'd130;
	sample_rom[239][20] = 8'd137;
	sample_rom[239][21] = 8'd139;
	sample_rom[239][22] = 8'd129;
	sample_rom[239][23] = 8'd119;
	sample_rom[239][24] = 8'd117;
	sample_rom[239][25] = 8'd121;
	sample_rom[239][26] = 8'd125;
	sample_rom[239][27] = 8'd128;
	sample_rom[239][28] = 8'd133;
	sample_rom[239][29] = 8'd138;
	sample_rom[239][30] = 8'd144;
	sample_rom[239][31] = 8'd136;
	sample_rom[239][32] = 8'd129;
	sample_rom[239][33] = 8'd126;
	sample_rom[239][34] = 8'd126;
	sample_rom[239][35] = 8'd128;
	sample_rom[239][36] = 8'd128;
	sample_rom[239][37] = 8'd128;
	sample_rom[239][38] = 8'd128;
	sample_rom[239][39] = 8'd133;
	sample_rom[239][40] = 8'd130;
	sample_rom[239][41] = 8'd127;
	sample_rom[239][42] = 8'd124;
	sample_rom[239][43] = 8'd124;
	sample_rom[239][44] = 8'd127;
	sample_rom[239][45] = 8'd124;
	sample_rom[239][46] = 8'd120;
	sample_rom[239][47] = 8'd123;
	sample_rom[239][48] = 8'd126;
	sample_rom[239][49] = 8'd129;
	sample_rom[239][50] = 8'd127;
	sample_rom[239][51] = 8'd127;
	sample_rom[239][52] = 8'd129;
	sample_rom[239][53] = 8'd134;
	sample_rom[239][54] = 8'd132;
	sample_rom[239][55] = 8'd131;
	sample_rom[239][56] = 8'd126;
	sample_rom[239][57] = 8'd128;
	sample_rom[239][58] = 8'd130;
	sample_rom[239][59] = 8'd132;
	sample_rom[239][60] = 8'd128;
	sample_rom[239][61] = 8'd131;
	sample_rom[239][62] = 8'd132;
	sample_rom[239][63] = 8'd134;
	sample_rom[240][0] = 8'd128;
	sample_rom[240][1] = 8'd207;
	sample_rom[240][2] = 8'd203;
	sample_rom[240][3] = 8'd132;
	sample_rom[240][4] = 8'd82;
	sample_rom[240][5] = 8'd97;
	sample_rom[240][6] = 8'd138;
	sample_rom[240][7] = 8'd146;
	sample_rom[240][8] = 8'd120;
	sample_rom[240][9] = 8'd110;
	sample_rom[240][10] = 8'd135;
	sample_rom[240][11] = 8'd162;
	sample_rom[240][12] = 8'd161;
	sample_rom[240][13] = 8'd133;
	sample_rom[240][14] = 8'd108;
	sample_rom[240][15] = 8'd106;
	sample_rom[240][16] = 8'd116;
	sample_rom[240][17] = 8'd122;
	sample_rom[240][18] = 8'd124;
	sample_rom[240][19] = 8'd130;
	sample_rom[240][20] = 8'd137;
	sample_rom[240][21] = 8'd139;
	sample_rom[240][22] = 8'd129;
	sample_rom[240][23] = 8'd119;
	sample_rom[240][24] = 8'd117;
	sample_rom[240][25] = 8'd121;
	sample_rom[240][26] = 8'd125;
	sample_rom[240][27] = 8'd128;
	sample_rom[240][28] = 8'd133;
	sample_rom[240][29] = 8'd138;
	sample_rom[240][30] = 8'd144;
	sample_rom[240][31] = 8'd136;
	sample_rom[240][32] = 8'd129;
	sample_rom[240][33] = 8'd126;
	sample_rom[240][34] = 8'd126;
	sample_rom[240][35] = 8'd128;
	sample_rom[240][36] = 8'd128;
	sample_rom[240][37] = 8'd128;
	sample_rom[240][38] = 8'd128;
	sample_rom[240][39] = 8'd133;
	sample_rom[240][40] = 8'd130;
	sample_rom[240][41] = 8'd127;
	sample_rom[240][42] = 8'd124;
	sample_rom[240][43] = 8'd124;
	sample_rom[240][44] = 8'd127;
	sample_rom[240][45] = 8'd124;
	sample_rom[240][46] = 8'd120;
	sample_rom[240][47] = 8'd123;
	sample_rom[240][48] = 8'd126;
	sample_rom[240][49] = 8'd129;
	sample_rom[240][50] = 8'd127;
	sample_rom[240][51] = 8'd127;
	sample_rom[240][52] = 8'd129;
	sample_rom[240][53] = 8'd134;
	sample_rom[240][54] = 8'd132;
	sample_rom[240][55] = 8'd131;
	sample_rom[240][56] = 8'd126;
	sample_rom[240][57] = 8'd128;
	sample_rom[240][58] = 8'd130;
	sample_rom[240][59] = 8'd132;
	sample_rom[240][60] = 8'd128;
	sample_rom[240][61] = 8'd131;
	sample_rom[240][62] = 8'd132;
	sample_rom[240][63] = 8'd134;
	sample_rom[241][0] = 8'd26;
	sample_rom[241][1] = 8'd16;
	sample_rom[241][2] = 8'd16;
	sample_rom[241][3] = 8'd206;
	sample_rom[241][4] = 8'd2;
	sample_rom[241][5] = 8'd0;
	sample_rom[241][6] = 8'd150;
	sample_rom[241][7] = 8'd8;
	sample_rom[241][8] = 8'd142;
	sample_rom[241][9] = 8'd3;
	sample_rom[241][10] = 8'd255;
	sample_rom[241][11] = 8'd111;
	sample_rom[241][12] = 8'd132;
	sample_rom[241][13] = 8'd48;
	sample_rom[241][14] = 8'd31;
	sample_rom[241][15] = 8'd38;
	sample_rom[241][16] = 8'd250;
	sample_rom[241][17] = 8'd111;
	sample_rom[241][18] = 8'd132;
	sample_rom[241][19] = 8'd151;
	sample_rom[241][20] = 8'd8;
	sample_rom[241][21] = 8'd189;
	sample_rom[241][22] = 8'd193;
	sample_rom[241][23] = 8'd66;
	sample_rom[241][24] = 8'd127;
	sample_rom[241][25] = 8'd176;
	sample_rom[241][26] = 8'd43;
	sample_rom[241][27] = 8'd127;
	sample_rom[241][28] = 8'd176;
	sample_rom[241][29] = 8'd42;
	sample_rom[241][30] = 8'd134;
	sample_rom[241][31] = 8'd4;
	sample_rom[241][32] = 8'd183;
	sample_rom[241][33] = 8'd176;
	sample_rom[241][34] = 8'd43;
	sample_rom[241][35] = 8'd141;
	sample_rom[241][36] = 8'd75;
	sample_rom[241][37] = 8'd134;
	sample_rom[241][38] = 8'd223;
	sample_rom[241][39] = 8'd183;
	sample_rom[241][40] = 8'd176;
	sample_rom[241][41] = 8'd113;
	sample_rom[241][42] = 8'd134;
	sample_rom[241][43] = 8'd255;
	sample_rom[241][44] = 8'd183;
	sample_rom[241][45] = 8'd2;
	sample_rom[241][46] = 8'd41;
	sample_rom[241][47] = 8'd134;
	sample_rom[241][48] = 8'd99;
	sample_rom[241][49] = 8'd151;
	sample_rom[241][50] = 8'd20;
	sample_rom[241][51] = 8'd134;
	sample_rom[241][52] = 8'd30;
	sample_rom[241][53] = 8'd138;
	sample_rom[241][54] = 8'd128;
	sample_rom[241][55] = 8'd151;
	sample_rom[241][56] = 8'd66;
	sample_rom[241][57] = 8'd182;
	sample_rom[241][58] = 8'd176;
	sample_rom[241][59] = 8'd112;
	sample_rom[241][60] = 8'd133;
	sample_rom[241][61] = 8'd4;
	sample_rom[241][62] = 8'd39;
	sample_rom[241][63] = 8'd6;
	sample_rom[242][0] = 8'd127;
	sample_rom[242][1] = 8'd60;
	sample_rom[242][2] = 8'd12;
	sample_rom[242][3] = 8'd124;
	sample_rom[242][4] = 8'd2;
	sample_rom[242][5] = 8'd107;
	sample_rom[242][6] = 8'd189;
	sample_rom[242][7] = 8'd215;
	sample_rom[242][8] = 8'd3;
	sample_rom[242][9] = 8'd189;
	sample_rom[242][10] = 8'd207;
	sample_rom[242][11] = 8'd0;
	sample_rom[242][12] = 8'd189;
	sample_rom[242][13] = 8'd196;
	sample_rom[242][14] = 8'd0;
	sample_rom[242][15] = 8'd189;
	sample_rom[242][16] = 8'd225;
	sample_rom[242][17] = 8'd21;
	sample_rom[242][18] = 8'd189;
	sample_rom[242][19] = 8'd174;
	sample_rom[242][20] = 8'd0;
	sample_rom[242][21] = 8'd150;
	sample_rom[242][22] = 8'd67;
	sample_rom[242][23] = 8'd133;
	sample_rom[242][24] = 8'd128;
	sample_rom[242][25] = 8'd39;
	sample_rom[242][26] = 8'd10;
	sample_rom[242][27] = 8'd150;
	sample_rom[242][28] = 8'd46;
	sample_rom[242][29] = 8'd52;
	sample_rom[242][30] = 8'd2;
	sample_rom[242][31] = 8'd141;
	sample_rom[242][32] = 8'd67;
	sample_rom[242][33] = 8'd53;
	sample_rom[242][34] = 8'd2;
	sample_rom[242][35] = 8'd151;
	sample_rom[242][36] = 8'd46;
	sample_rom[242][37] = 8'd189;
	sample_rom[242][38] = 8'd236;
	sample_rom[242][39] = 8'd0;
	sample_rom[242][40] = 8'd189;
	sample_rom[242][41] = 8'd208;
	sample_rom[242][42] = 8'd0;
	sample_rom[242][43] = 8'd189;
	sample_rom[242][44] = 8'd210;
	sample_rom[242][45] = 8'd0;
	sample_rom[242][46] = 8'd32;
	sample_rom[242][47] = 8'd214;
	sample_rom[242][48] = 8'd26;
	sample_rom[242][49] = 8'd16;
	sample_rom[242][50] = 8'd190;
	sample_rom[242][51] = 8'd239;
	sample_rom[242][52] = 8'd248;
	sample_rom[242][53] = 8'd191;
	sample_rom[242][54] = 8'd191;
	sample_rom[242][55] = 8'd150;
	sample_rom[242][56] = 8'd134;
	sample_rom[242][57] = 8'd129;
	sample_rom[242][58] = 8'd183;
	sample_rom[242][59] = 8'd176;
	sample_rom[242][60] = 8'd81;
	sample_rom[242][61] = 8'd198;
	sample_rom[242][62] = 8'd208;
	sample_rom[242][63] = 8'd247;
	sample_rom[243][0] = 8'd176;
	sample_rom[243][1] = 8'd80;
	sample_rom[243][2] = 8'd134;
	sample_rom[243][3] = 8'd128;
	sample_rom[243][4] = 8'd183;
	sample_rom[243][5] = 8'd176;
	sample_rom[243][6] = 8'd81;
	sample_rom[243][7] = 8'd198;
	sample_rom[243][8] = 8'd146;
	sample_rom[243][9] = 8'd247;
	sample_rom[243][10] = 8'd176;
	sample_rom[243][11] = 8'd80;
	sample_rom[243][12] = 8'd134;
	sample_rom[243][13] = 8'd160;
	sample_rom[243][14] = 8'd183;
	sample_rom[243][15] = 8'd176;
	sample_rom[243][16] = 8'd126;
	sample_rom[243][17] = 8'd134;
	sample_rom[243][18] = 8'd113;
	sample_rom[243][19] = 8'd183;
	sample_rom[243][20] = 8'd176;
	sample_rom[243][21] = 8'd114;
	sample_rom[243][22] = 8'd134;
	sample_rom[243][23] = 8'd128;
	sample_rom[243][24] = 8'd183;
	sample_rom[243][25] = 8'd176;
	sample_rom[243][26] = 8'd112;
	sample_rom[243][27] = 8'd134;
	sample_rom[243][28] = 8'd0;
	sample_rom[243][29] = 8'd183;
	sample_rom[243][30] = 8'd176;
	sample_rom[243][31] = 8'd37;
	sample_rom[243][32] = 8'd141;
	sample_rom[243][33] = 8'd2;
	sample_rom[243][34] = 8'd32;
	sample_rom[243][35] = 8'd45;
	sample_rom[243][36] = 8'd79;
	sample_rom[243][37] = 8'd142;
	sample_rom[243][38] = 8'd0;
	sample_rom[243][39] = 8'd224;
	sample_rom[243][40] = 8'd141;
	sample_rom[243][41] = 8'd27;
	sample_rom[243][42] = 8'd142;
	sample_rom[243][43] = 8'd0;
	sample_rom[243][44] = 8'd136;
	sample_rom[243][45] = 8'd141;
	sample_rom[243][46] = 8'd22;
	sample_rom[243][47] = 8'd142;
	sample_rom[243][48] = 8'd0;
	sample_rom[243][49] = 8'd248;
	sample_rom[243][50] = 8'd141;
	sample_rom[243][51] = 8'd17;
	sample_rom[243][52] = 8'd134;
	sample_rom[243][53] = 8'd64;
	sample_rom[243][54] = 8'd142;
	sample_rom[243][55] = 8'd0;
	sample_rom[243][56] = 8'd152;
	sample_rom[243][57] = 8'd141;
	sample_rom[243][58] = 8'd10;
	sample_rom[243][59] = 8'd142;
	sample_rom[243][60] = 8'd0;
	sample_rom[243][61] = 8'd232;
	sample_rom[243][62] = 8'd141;
	sample_rom[243][63] = 8'd5;
	sample_rom[244][0] = 8'd122;
	sample_rom[244][1] = 8'd121;
	sample_rom[244][2] = 8'd121;
	sample_rom[244][3] = 8'd122;
	sample_rom[244][4] = 8'd123;
	sample_rom[244][5] = 8'd123;
	sample_rom[244][6] = 8'd123;
	sample_rom[244][7] = 8'd124;
	sample_rom[244][8] = 8'd124;
	sample_rom[244][9] = 8'd125;
	sample_rom[244][10] = 8'd125;
	sample_rom[244][11] = 8'd125;
	sample_rom[244][12] = 8'd125;
	sample_rom[244][13] = 8'd126;
	sample_rom[244][14] = 8'd126;
	sample_rom[244][15] = 8'd126;
	sample_rom[244][16] = 8'd126;
	sample_rom[244][17] = 8'd125;
	sample_rom[244][18] = 8'd126;
	sample_rom[244][19] = 8'd126;
	sample_rom[244][20] = 8'd127;
	sample_rom[244][21] = 8'd127;
	sample_rom[244][22] = 8'd127;
	sample_rom[244][23] = 8'd127;
	sample_rom[244][24] = 8'd127;
	sample_rom[244][25] = 8'd126;
	sample_rom[244][26] = 8'd125;
	sample_rom[244][27] = 8'd125;
	sample_rom[244][28] = 8'd124;
	sample_rom[244][29] = 8'd124;
	sample_rom[244][30] = 8'd123;
	sample_rom[244][31] = 8'd123;
	sample_rom[244][32] = 8'd123;
	sample_rom[244][33] = 8'd123;
	sample_rom[244][34] = 8'd124;
	sample_rom[244][35] = 8'd124;
	sample_rom[244][36] = 8'd125;
	sample_rom[244][37] = 8'd125;
	sample_rom[244][38] = 8'd125;
	sample_rom[244][39] = 8'd125;
	sample_rom[244][40] = 8'd125;
	sample_rom[244][41] = 8'd124;
	sample_rom[244][42] = 8'd123;
	sample_rom[244][43] = 8'd125;
	sample_rom[244][44] = 8'd125;
	sample_rom[244][45] = 8'd120;
	sample_rom[244][46] = 8'd119;
	sample_rom[244][47] = 8'd123;
	sample_rom[244][48] = 8'd125;
	sample_rom[244][49] = 8'd121;
	sample_rom[244][50] = 8'd119;
	sample_rom[244][51] = 8'd124;
	sample_rom[244][52] = 8'd127;
	sample_rom[244][53] = 8'd118;
	sample_rom[244][54] = 8'd113;
	sample_rom[244][55] = 8'd119;
	sample_rom[244][56] = 8'd125;
	sample_rom[244][57] = 8'd117;
	sample_rom[244][58] = 8'd104;
	sample_rom[244][59] = 8'd113;
	sample_rom[244][60] = 8'd120;
	sample_rom[244][61] = 8'd119;
	sample_rom[244][62] = 8'd117;
	sample_rom[244][63] = 8'd119;
	sample_rom[245][0] = 8'd115;
	sample_rom[245][1] = 8'd101;
	sample_rom[245][2] = 8'd94;
	sample_rom[245][3] = 8'd86;
	sample_rom[245][4] = 8'd91;
	sample_rom[245][5] = 8'd109;
	sample_rom[245][6] = 8'd120;
	sample_rom[245][7] = 8'd129;
	sample_rom[245][8] = 8'd130;
	sample_rom[245][9] = 8'd121;
	sample_rom[245][10] = 8'd131;
	sample_rom[245][11] = 8'd148;
	sample_rom[245][12] = 8'd150;
	sample_rom[245][13] = 8'd141;
	sample_rom[245][14] = 8'd131;
	sample_rom[245][15] = 8'd136;
	sample_rom[245][16] = 8'd169;
	sample_rom[245][17] = 8'd181;
	sample_rom[245][18] = 8'd160;
	sample_rom[245][19] = 8'd134;
	sample_rom[245][20] = 8'd123;
	sample_rom[245][21] = 8'd103;
	sample_rom[245][22] = 8'd84;
	sample_rom[245][23] = 8'd71;
	sample_rom[245][24] = 8'd75;
	sample_rom[245][25] = 8'd72;
	sample_rom[245][26] = 8'd84;
	sample_rom[245][27] = 8'd104;
	sample_rom[245][28] = 8'd108;
	sample_rom[245][29] = 8'd107;
	sample_rom[245][30] = 8'd134;
	sample_rom[245][31] = 8'd181;
	sample_rom[245][32] = 8'd197;
	sample_rom[245][33] = 8'd183;
	sample_rom[245][34] = 8'd184;
	sample_rom[245][35] = 8'd204;
	sample_rom[245][36] = 8'd212;
	sample_rom[245][37] = 8'd203;
	sample_rom[245][38] = 8'd201;
	sample_rom[245][39] = 8'd186;
	sample_rom[245][40] = 8'd161;
	sample_rom[245][41] = 8'd155;
	sample_rom[245][42] = 8'd169;
	sample_rom[245][43] = 8'd168;
	sample_rom[245][44] = 8'd151;
	sample_rom[245][45] = 8'd120;
	sample_rom[245][46] = 8'd106;
	sample_rom[245][47] = 8'd97;
	sample_rom[245][48] = 8'd100;
	sample_rom[245][49] = 8'd84;
	sample_rom[245][50] = 8'd74;
	sample_rom[245][51] = 8'd96;
	sample_rom[245][52] = 8'd111;
	sample_rom[245][53] = 8'd117;
	sample_rom[245][54] = 8'd104;
	sample_rom[245][55] = 8'd90;
	sample_rom[245][56] = 8'd63;
	sample_rom[245][57] = 8'd46;
	sample_rom[245][58] = 8'd52;
	sample_rom[245][59] = 8'd73;
	sample_rom[245][60] = 8'd79;
	sample_rom[245][61] = 8'd65;
	sample_rom[245][62] = 8'd45;
	sample_rom[245][63] = 8'd37;
	sample_rom[246][0] = 8'd24;
	sample_rom[246][1] = 8'd14;
	sample_rom[246][2] = 8'd23;
	sample_rom[246][3] = 8'd8;
	sample_rom[246][4] = 8'd7;
	sample_rom[246][5] = 8'd43;
	sample_rom[246][6] = 8'd73;
	sample_rom[246][7] = 8'd76;
	sample_rom[246][8] = 8'd62;
	sample_rom[246][9] = 8'd77;
	sample_rom[246][10] = 8'd110;
	sample_rom[246][11] = 8'd141;
	sample_rom[246][12] = 8'd168;
	sample_rom[246][13] = 8'd189;
	sample_rom[246][14] = 8'd213;
	sample_rom[246][15] = 8'd222;
	sample_rom[246][16] = 8'd218;
	sample_rom[246][17] = 8'd226;
	sample_rom[246][18] = 8'd225;
	sample_rom[246][19] = 8'd225;
	sample_rom[246][20] = 8'd223;
	sample_rom[246][21] = 8'd223;
	sample_rom[246][22] = 8'd212;
	sample_rom[246][23] = 8'd164;
	sample_rom[246][24] = 8'd134;
	sample_rom[246][25] = 8'd147;
	sample_rom[246][26] = 8'd156;
	sample_rom[246][27] = 8'd133;
	sample_rom[246][28] = 8'd97;
	sample_rom[246][29] = 8'd91;
	sample_rom[246][30] = 8'd118;
	sample_rom[246][31] = 8'd122;
	sample_rom[246][32] = 8'd106;
	sample_rom[246][33] = 8'd84;
	sample_rom[246][34] = 8'd75;
	sample_rom[246][35] = 8'd103;
	sample_rom[246][36] = 8'd145;
	sample_rom[246][37] = 8'd188;
	sample_rom[246][38] = 8'd192;
	sample_rom[246][39] = 8'd160;
	sample_rom[246][40] = 8'd152;
	sample_rom[246][41] = 8'd166;
	sample_rom[246][42] = 8'd198;
	sample_rom[246][43] = 8'd203;
	sample_rom[246][44] = 8'd197;
	sample_rom[246][45] = 8'd181;
	sample_rom[246][46] = 8'd145;
	sample_rom[246][47] = 8'd120;
	sample_rom[246][48] = 8'd118;
	sample_rom[246][49] = 8'd126;
	sample_rom[246][50] = 8'd130;
	sample_rom[246][51] = 8'd141;
	sample_rom[246][52] = 8'd162;
	sample_rom[246][53] = 8'd139;
	sample_rom[246][54] = 8'd89;
	sample_rom[246][55] = 8'd53;
	sample_rom[246][56] = 8'd45;
	sample_rom[246][57] = 8'd49;
	sample_rom[246][58] = 8'd35;
	sample_rom[246][59] = 8'd23;
	sample_rom[246][60] = 8'd49;
	sample_rom[246][61] = 8'd42;
	sample_rom[246][62] = 8'd4;
	sample_rom[246][63] = 8'd0;
	sample_rom[247][0] = 8'd0;
	sample_rom[247][1] = 8'd0;
	sample_rom[247][2] = 8'd0;
	sample_rom[247][3] = 8'd0;
	sample_rom[247][4] = 8'd19;
	sample_rom[247][5] = 8'd62;
	sample_rom[247][6] = 8'd53;
	sample_rom[247][7] = 8'd21;
	sample_rom[247][8] = 8'd31;
	sample_rom[247][9] = 8'd70;
	sample_rom[247][10] = 8'd121;
	sample_rom[247][11] = 8'd172;
	sample_rom[247][12] = 8'd219;
	sample_rom[247][13] = 8'd228;
	sample_rom[247][14] = 8'd228;
	sample_rom[247][15] = 8'd227;
	sample_rom[247][16] = 8'd220;
	sample_rom[247][17] = 8'd223;
	sample_rom[247][18] = 8'd225;
	sample_rom[247][19] = 8'd224;
	sample_rom[247][20] = 8'd223;
	sample_rom[247][21] = 8'd218;
	sample_rom[247][22] = 8'd190;
	sample_rom[247][23] = 8'd140;
	sample_rom[247][24] = 8'd89;
	sample_rom[247][25] = 8'd62;
	sample_rom[247][26] = 8'd71;
	sample_rom[247][27] = 8'd69;
	sample_rom[247][28] = 8'd50;
	sample_rom[247][29] = 8'd51;
	sample_rom[247][30] = 8'd73;
	sample_rom[247][31] = 8'd83;
	sample_rom[247][32] = 8'd40;
	sample_rom[247][33] = 8'd1;
	sample_rom[247][34] = 8'd29;
	sample_rom[247][35] = 8'd103;
	sample_rom[247][36] = 8'd183;
	sample_rom[247][37] = 8'd201;
	sample_rom[247][38] = 8'd198;
	sample_rom[247][39] = 8'd219;
	sample_rom[247][40] = 8'd224;
	sample_rom[247][41] = 8'd224;
	sample_rom[247][42] = 8'd222;
	sample_rom[247][43] = 8'd221;
	sample_rom[247][44] = 8'd221;
	sample_rom[247][45] = 8'd220;
	sample_rom[247][46] = 8'd212;
	sample_rom[247][47] = 8'd191;
	sample_rom[247][48] = 8'd168;
	sample_rom[247][49] = 8'd144;
	sample_rom[247][50] = 8'd129;
	sample_rom[247][51] = 8'd155;
	sample_rom[247][52] = 8'd178;
	sample_rom[247][53] = 8'd143;
	sample_rom[247][54] = 8'd89;
	sample_rom[247][55] = 8'd57;
	sample_rom[247][56] = 8'd50;
	sample_rom[247][57] = 8'd46;
	sample_rom[247][58] = 8'd45;
	sample_rom[247][59] = 8'd53;
	sample_rom[247][60] = 8'd47;
	sample_rom[247][61] = 8'd28;
	sample_rom[247][62] = 8'd6;
	sample_rom[247][63] = 8'd0;
	sample_rom[248][0] = 8'd0;
	sample_rom[248][1] = 8'd0;
	sample_rom[248][2] = 8'd0;
	sample_rom[248][3] = 8'd0;
	sample_rom[248][4] = 8'd24;
	sample_rom[248][5] = 8'd51;
	sample_rom[248][6] = 8'd48;
	sample_rom[248][7] = 8'd39;
	sample_rom[248][8] = 8'd58;
	sample_rom[248][9] = 8'd98;
	sample_rom[248][10] = 8'd145;
	sample_rom[248][11] = 8'd185;
	sample_rom[248][12] = 8'd215;
	sample_rom[248][13] = 8'd230;
	sample_rom[248][14] = 8'd229;
	sample_rom[248][15] = 8'd217;
	sample_rom[248][16] = 8'd201;
	sample_rom[248][17] = 8'd223;
	sample_rom[248][18] = 8'd226;
	sample_rom[248][19] = 8'd225;
	sample_rom[248][20] = 8'd224;
	sample_rom[248][21] = 8'd211;
	sample_rom[248][22] = 8'd181;
	sample_rom[248][23] = 8'd139;
	sample_rom[248][24] = 8'd86;
	sample_rom[248][25] = 8'd64;
	sample_rom[248][26] = 8'd61;
	sample_rom[248][27] = 8'd47;
	sample_rom[248][28] = 8'd45;
	sample_rom[248][29] = 8'd61;
	sample_rom[248][30] = 8'd91;
	sample_rom[248][31] = 8'd77;
	sample_rom[248][32] = 8'd24;
	sample_rom[248][33] = 8'd29;
	sample_rom[248][34] = 8'd99;
	sample_rom[248][35] = 8'd169;
	sample_rom[248][36] = 8'd184;
	sample_rom[248][37] = 8'd187;
	sample_rom[248][38] = 8'd220;
	sample_rom[248][39] = 8'd225;
	sample_rom[248][40] = 8'd225;
	sample_rom[248][41] = 8'd224;
	sample_rom[248][42] = 8'd223;
	sample_rom[248][43] = 8'd222;
	sample_rom[248][44] = 8'd222;
	sample_rom[248][45] = 8'd216;
	sample_rom[248][46] = 8'd187;
	sample_rom[248][47] = 8'd163;
	sample_rom[248][48] = 8'd147;
	sample_rom[248][49] = 8'd146;
	sample_rom[248][50] = 8'd162;
	sample_rom[248][51] = 8'd170;
	sample_rom[248][52] = 8'd162;
	sample_rom[248][53] = 8'd136;
	sample_rom[248][54] = 8'd96;
	sample_rom[248][55] = 8'd64;
	sample_rom[248][56] = 8'd76;
	sample_rom[248][57] = 8'd99;
	sample_rom[248][58] = 8'd102;
	sample_rom[248][59] = 8'd88;
	sample_rom[248][60] = 8'd80;
	sample_rom[248][61] = 8'd72;
	sample_rom[248][62] = 8'd42;
	sample_rom[248][63] = 8'd7;
	sample_rom[249][0] = 8'd0;
	sample_rom[249][1] = 8'd0;
	sample_rom[249][2] = 8'd0;
	sample_rom[249][3] = 8'd0;
	sample_rom[249][4] = 8'd27;
	sample_rom[249][5] = 8'd30;
	sample_rom[249][6] = 8'd5;
	sample_rom[249][7] = 8'd2;
	sample_rom[249][8] = 8'd23;
	sample_rom[249][9] = 8'd55;
	sample_rom[249][10] = 8'd93;
	sample_rom[249][11] = 8'd141;
	sample_rom[249][12] = 8'd199;
	sample_rom[249][13] = 8'd214;
	sample_rom[249][14] = 8'd197;
	sample_rom[249][15] = 8'd182;
	sample_rom[249][16] = 8'd209;
	sample_rom[249][17] = 8'd228;
	sample_rom[249][18] = 8'd227;
	sample_rom[249][19] = 8'd227;
	sample_rom[249][20] = 8'd225;
	sample_rom[249][21] = 8'd224;
	sample_rom[249][22] = 8'd209;
	sample_rom[249][23] = 8'd166;
	sample_rom[249][24] = 8'd128;
	sample_rom[249][25] = 8'd102;
	sample_rom[249][26] = 8'd70;
	sample_rom[249][27] = 8'd60;
	sample_rom[249][28] = 8'd82;
	sample_rom[249][29] = 8'd115;
	sample_rom[249][30] = 8'd83;
	sample_rom[249][31] = 8'd24;
	sample_rom[249][32] = 8'd8;
	sample_rom[249][33] = 8'd39;
	sample_rom[249][34] = 8'd79;
	sample_rom[249][35] = 8'd107;
	sample_rom[249][36] = 8'd117;
	sample_rom[249][37] = 8'd147;
	sample_rom[249][38] = 8'd172;
	sample_rom[249][39] = 8'd182;
	sample_rom[249][40] = 8'd188;
	sample_rom[249][41] = 8'd213;
	sample_rom[249][42] = 8'd225;
	sample_rom[249][43] = 8'd224;
	sample_rom[249][44] = 8'd224;
	sample_rom[249][45] = 8'd208;
	sample_rom[249][46] = 8'd175;
	sample_rom[249][47] = 8'd173;
	sample_rom[249][48] = 8'd186;
	sample_rom[249][49] = 8'd183;
	sample_rom[249][50] = 8'd187;
	sample_rom[249][51] = 8'd201;
	sample_rom[249][52] = 8'd197;
	sample_rom[249][53] = 8'd155;
	sample_rom[249][54] = 8'd109;
	sample_rom[249][55] = 8'd111;
	sample_rom[249][56] = 8'd130;
	sample_rom[249][57] = 8'd128;
	sample_rom[249][58] = 8'd112;
	sample_rom[249][59] = 8'd104;
	sample_rom[249][60] = 8'd105;
	sample_rom[249][61] = 8'd72;
	sample_rom[249][62] = 8'd23;
	sample_rom[249][63] = 8'd0;
	sample_rom[250][0] = 8'd0;
	sample_rom[250][1] = 8'd0;
	sample_rom[250][2] = 8'd0;
	sample_rom[250][3] = 8'd3;
	sample_rom[250][4] = 8'd9;
	sample_rom[250][5] = 8'd0;
	sample_rom[250][6] = 8'd0;
	sample_rom[250][7] = 8'd0;
	sample_rom[250][8] = 8'd7;
	sample_rom[250][9] = 8'd38;
	sample_rom[250][10] = 8'd85;
	sample_rom[250][11] = 8'd142;
	sample_rom[250][12] = 8'd180;
	sample_rom[250][13] = 8'd190;
	sample_rom[250][14] = 8'd190;
	sample_rom[250][15] = 8'd205;
	sample_rom[250][16] = 8'd228;
	sample_rom[250][17] = 8'd228;
	sample_rom[250][18] = 8'd227;
	sample_rom[250][19] = 8'd227;
	sample_rom[250][20] = 8'd225;
	sample_rom[250][21] = 8'd225;
	sample_rom[250][22] = 8'd224;
	sample_rom[250][23] = 8'd192;
	sample_rom[250][24] = 8'd140;
	sample_rom[250][25] = 8'd79;
	sample_rom[250][26] = 8'd68;
	sample_rom[250][27] = 8'd102;
	sample_rom[250][28] = 8'd112;
	sample_rom[250][29] = 8'd84;
	sample_rom[250][30] = 8'd40;
	sample_rom[250][31] = 8'd18;
	sample_rom[250][32] = 8'd21;
	sample_rom[250][33] = 8'd42;
	sample_rom[250][34] = 8'd73;
	sample_rom[250][35] = 8'd107;
	sample_rom[250][36] = 8'd127;
	sample_rom[250][37] = 8'd137;
	sample_rom[250][38] = 8'd162;
	sample_rom[250][39] = 8'd185;
	sample_rom[250][40] = 8'd191;
	sample_rom[250][41] = 8'd202;
	sample_rom[250][42] = 8'd225;
	sample_rom[250][43] = 8'd225;
	sample_rom[250][44] = 8'd210;
	sample_rom[250][45] = 8'd172;
	sample_rom[250][46] = 8'd168;
	sample_rom[250][47] = 8'd172;
	sample_rom[250][48] = 8'd154;
	sample_rom[250][49] = 8'd153;
	sample_rom[250][50] = 8'd172;
	sample_rom[250][51] = 8'd178;
	sample_rom[250][52] = 8'd147;
	sample_rom[250][53] = 8'd100;
	sample_rom[250][54] = 8'd89;
	sample_rom[250][55] = 8'd99;
	sample_rom[250][56] = 8'd102;
	sample_rom[250][57] = 8'd101;
	sample_rom[250][58] = 8'd92;
	sample_rom[250][59] = 8'd106;
	sample_rom[250][60] = 8'd109;
	sample_rom[250][61] = 8'd80;
	sample_rom[250][62] = 8'd23;
	sample_rom[250][63] = 8'd0;
	sample_rom[251][0] = 8'd0;
	sample_rom[251][1] = 8'd0;
	sample_rom[251][2] = 8'd3;
	sample_rom[251][3] = 8'd15;
	sample_rom[251][4] = 8'd17;
	sample_rom[251][5] = 8'd9;
	sample_rom[251][6] = 8'd2;
	sample_rom[251][7] = 8'd0;
	sample_rom[251][8] = 8'd13;
	sample_rom[251][9] = 8'd60;
	sample_rom[251][10] = 8'd108;
	sample_rom[251][11] = 8'd139;
	sample_rom[251][12] = 8'd162;
	sample_rom[251][13] = 8'd179;
	sample_rom[251][14] = 8'd185;
	sample_rom[251][15] = 8'd211;
	sample_rom[251][16] = 8'd230;
	sample_rom[251][17] = 8'd230;
	sample_rom[251][18] = 8'd229;
	sample_rom[251][19] = 8'd229;
	sample_rom[251][20] = 8'd228;
	sample_rom[251][21] = 8'd227;
	sample_rom[251][22] = 8'd226;
	sample_rom[251][23] = 8'd185;
	sample_rom[251][24] = 8'd118;
	sample_rom[251][25] = 8'd107;
	sample_rom[251][26] = 8'd143;
	sample_rom[251][27] = 8'd153;
	sample_rom[251][28] = 8'd127;
	sample_rom[251][29] = 8'd96;
	sample_rom[251][30] = 8'd78;
	sample_rom[251][31] = 8'd57;
	sample_rom[251][32] = 8'd43;
	sample_rom[251][33] = 8'd67;
	sample_rom[251][34] = 8'd106;
	sample_rom[251][35] = 8'd119;
	sample_rom[251][36] = 8'd128;
	sample_rom[251][37] = 8'd154;
	sample_rom[251][38] = 8'd178;
	sample_rom[251][39] = 8'd179;
	sample_rom[251][40] = 8'd186;
	sample_rom[251][41] = 8'd220;
	sample_rom[251][42] = 8'd226;
	sample_rom[251][43] = 8'd219;
	sample_rom[251][44] = 8'd190;
	sample_rom[251][45] = 8'd160;
	sample_rom[251][46] = 8'd151;
	sample_rom[251][47] = 8'd139;
	sample_rom[251][48] = 8'd140;
	sample_rom[251][49] = 8'd151;
	sample_rom[251][50] = 8'd157;
	sample_rom[251][51] = 8'd152;
	sample_rom[251][52] = 8'd117;
	sample_rom[251][53] = 8'd91;
	sample_rom[251][54] = 8'd88;
	sample_rom[251][55] = 8'd105;
	sample_rom[251][56] = 8'd108;
	sample_rom[251][57] = 8'd96;
	sample_rom[251][58] = 8'd112;
	sample_rom[251][59] = 8'd138;
	sample_rom[251][60] = 8'd127;
	sample_rom[251][61] = 8'd72;
	sample_rom[251][62] = 8'd23;
	sample_rom[251][63] = 8'd11;
	sample_rom[252][0] = 8'd17;
	sample_rom[252][1] = 8'd15;
	sample_rom[252][2] = 8'd19;
	sample_rom[252][3] = 8'd35;
	sample_rom[252][4] = 8'd41;
	sample_rom[252][5] = 8'd14;
	sample_rom[252][6] = 8'd0;
	sample_rom[252][7] = 8'd0;
	sample_rom[252][8] = 8'd19;
	sample_rom[252][9] = 8'd66;
	sample_rom[252][10] = 8'd97;
	sample_rom[252][11] = 8'd113;
	sample_rom[252][12] = 8'd142;
	sample_rom[252][13] = 8'd164;
	sample_rom[252][14] = 8'd169;
	sample_rom[252][15] = 8'd206;
	sample_rom[252][16] = 8'd230;
	sample_rom[252][17] = 8'd230;
	sample_rom[252][18] = 8'd230;
	sample_rom[252][19] = 8'd229;
	sample_rom[252][20] = 8'd228;
	sample_rom[252][21] = 8'd227;
	sample_rom[252][22] = 8'd226;
	sample_rom[252][23] = 8'd156;
	sample_rom[252][24] = 8'd127;
	sample_rom[252][25] = 8'd153;
	sample_rom[252][26] = 8'd163;
	sample_rom[252][27] = 8'd146;
	sample_rom[252][28] = 8'd129;
	sample_rom[252][29] = 8'd108;
	sample_rom[252][30] = 8'd80;
	sample_rom[252][31] = 8'd52;
	sample_rom[252][32] = 8'd53;
	sample_rom[252][33] = 8'd78;
	sample_rom[252][34] = 8'd96;
	sample_rom[252][35] = 8'd124;
	sample_rom[252][36] = 8'd135;
	sample_rom[252][37] = 8'd151;
	sample_rom[252][38] = 8'd167;
	sample_rom[252][39] = 8'd181;
	sample_rom[252][40] = 8'd202;
	sample_rom[252][41] = 8'd215;
	sample_rom[252][42] = 8'd225;
	sample_rom[252][43] = 8'd219;
	sample_rom[252][44] = 8'd188;
	sample_rom[252][45] = 8'd155;
	sample_rom[252][46] = 8'd148;
	sample_rom[252][47] = 8'd154;
	sample_rom[252][48] = 8'd155;
	sample_rom[252][49] = 8'd152;
	sample_rom[252][50] = 8'd155;
	sample_rom[252][51] = 8'd136;
	sample_rom[252][52] = 8'd105;
	sample_rom[252][53] = 8'd87;
	sample_rom[252][54] = 8'd82;
	sample_rom[252][55] = 8'd83;
	sample_rom[252][56] = 8'd79;
	sample_rom[252][57] = 8'd82;
	sample_rom[252][58] = 8'd103;
	sample_rom[252][59] = 8'd114;
	sample_rom[252][60] = 8'd84;
	sample_rom[252][61] = 8'd32;
	sample_rom[252][62] = 8'd9;
	sample_rom[252][63] = 8'd6;
	sample_rom[253][0] = 8'd6;
	sample_rom[253][1] = 8'd8;
	sample_rom[253][2] = 8'd27;
	sample_rom[253][3] = 8'd44;
	sample_rom[253][4] = 8'd38;
	sample_rom[253][5] = 8'd9;
	sample_rom[253][6] = 8'd0;
	sample_rom[253][7] = 8'd3;
	sample_rom[253][8] = 8'd44;
	sample_rom[253][9] = 8'd76;
	sample_rom[253][10] = 8'd104;
	sample_rom[253][11] = 8'd131;
	sample_rom[253][12] = 8'd146;
	sample_rom[253][13] = 8'd155;
	sample_rom[253][14] = 8'd191;
	sample_rom[253][15] = 8'd227;
	sample_rom[253][16] = 8'd233;
	sample_rom[253][17] = 8'd232;
	sample_rom[253][18] = 8'd232;
	sample_rom[253][19] = 8'd231;
	sample_rom[253][20] = 8'd229;
	sample_rom[253][21] = 8'd229;
	sample_rom[253][22] = 8'd206;
	sample_rom[253][23] = 8'd159;
	sample_rom[253][24] = 8'd152;
	sample_rom[253][25] = 8'd158;
	sample_rom[253][26] = 8'd161;
	sample_rom[253][27] = 8'd149;
	sample_rom[253][28] = 8'd115;
	sample_rom[253][29] = 8'd94;
	sample_rom[253][30] = 8'd73;
	sample_rom[253][31] = 8'd46;
	sample_rom[253][32] = 8'd38;
	sample_rom[253][33] = 8'd64;
	sample_rom[253][34] = 8'd102;
	sample_rom[253][35] = 8'd111;
	sample_rom[253][36] = 8'd113;
	sample_rom[253][37] = 8'd138;
	sample_rom[253][38] = 8'd166;
	sample_rom[253][39] = 8'd177;
	sample_rom[253][40] = 8'd188;
	sample_rom[253][41] = 8'd217;
	sample_rom[253][42] = 8'd226;
	sample_rom[253][43] = 8'd217;
	sample_rom[253][44] = 8'd185;
	sample_rom[253][45] = 8'd160;
	sample_rom[253][46] = 8'd165;
	sample_rom[253][47] = 8'd174;
	sample_rom[253][48] = 8'd168;
	sample_rom[253][49] = 8'd162;
	sample_rom[253][50] = 8'd161;
	sample_rom[253][51] = 8'd151;
	sample_rom[253][52] = 8'd127;
	sample_rom[253][53] = 8'd107;
	sample_rom[253][54] = 8'd98;
	sample_rom[253][55] = 8'd93;
	sample_rom[253][56] = 8'd94;
	sample_rom[253][57] = 8'd108;
	sample_rom[253][58] = 8'd119;
	sample_rom[253][59] = 8'd115;
	sample_rom[253][60] = 8'd78;
	sample_rom[253][61] = 8'd32;
	sample_rom[253][62] = 8'd9;
	sample_rom[253][63] = 8'd4;
	sample_rom[254][0] = 8'd2;
	sample_rom[254][1] = 8'd13;
	sample_rom[254][2] = 8'd42;
	sample_rom[254][3] = 8'd51;
	sample_rom[254][4] = 8'd23;
	sample_rom[254][5] = 8'd0;
	sample_rom[254][6] = 8'd0;
	sample_rom[254][7] = 8'd7;
	sample_rom[254][8] = 8'd50;
	sample_rom[254][9] = 8'd89;
	sample_rom[254][10] = 8'd103;
	sample_rom[254][11] = 8'd112;
	sample_rom[254][12] = 8'd132;
	sample_rom[254][13] = 8'd175;
	sample_rom[254][14] = 8'd213;
	sample_rom[254][15] = 8'd230;
	sample_rom[254][16] = 8'd232;
	sample_rom[254][17] = 8'd231;
	sample_rom[254][18] = 8'd230;
	sample_rom[254][19] = 8'd229;
	sample_rom[254][20] = 8'd228;
	sample_rom[254][21] = 8'd228;
	sample_rom[254][22] = 8'd190;
	sample_rom[254][23] = 8'd144;
	sample_rom[254][24] = 8'd148;
	sample_rom[254][25] = 8'd164;
	sample_rom[254][26] = 8'd151;
	sample_rom[254][27] = 8'd123;
	sample_rom[254][28] = 8'd111;
	sample_rom[254][29] = 8'd96;
	sample_rom[254][30] = 8'd55;
	sample_rom[254][31] = 8'd26;
	sample_rom[254][32] = 8'd41;
	sample_rom[254][33] = 8'd81;
	sample_rom[254][34] = 8'd94;
	sample_rom[254][35] = 8'd91;
	sample_rom[254][36] = 8'd113;
	sample_rom[254][37] = 8'd141;
	sample_rom[254][38] = 8'd159;
	sample_rom[254][39] = 8'd167;
	sample_rom[254][40] = 8'd192;
	sample_rom[254][41] = 8'd222;
	sample_rom[254][42] = 8'd226;
	sample_rom[254][43] = 8'd200;
	sample_rom[254][44] = 8'd167;
	sample_rom[254][45] = 8'd161;
	sample_rom[254][46] = 8'd174;
	sample_rom[254][47] = 8'd174;
	sample_rom[254][48] = 8'd162;
	sample_rom[254][49] = 8'd155;
	sample_rom[254][50] = 8'd157;
	sample_rom[254][51] = 8'd154;
	sample_rom[254][52] = 8'd123;
	sample_rom[254][53] = 8'd93;
	sample_rom[254][54] = 8'd86;
	sample_rom[254][55] = 8'd95;
	sample_rom[254][56] = 8'd101;
	sample_rom[254][57] = 8'd112;
	sample_rom[254][58] = 8'd119;
	sample_rom[254][59] = 8'd107;
	sample_rom[254][60] = 8'd75;
	sample_rom[254][61] = 8'd32;
	sample_rom[254][62] = 8'd8;
	sample_rom[254][63] = 8'd3;
	sample_rom[255][0] = 8'd21;
	sample_rom[255][1] = 8'd38;
	sample_rom[255][2] = 8'd53;
	sample_rom[255][3] = 8'd54;
	sample_rom[255][4] = 8'd27;
	sample_rom[255][5] = 8'd3;
	sample_rom[255][6] = 8'd0;
	sample_rom[255][7] = 8'd29;
	sample_rom[255][8] = 8'd80;
	sample_rom[255][9] = 8'd90;
	sample_rom[255][10] = 8'd80;
	sample_rom[255][11] = 8'd101;
	sample_rom[255][12] = 8'd156;
	sample_rom[255][13] = 8'd187;
	sample_rom[255][14] = 8'd190;
	sample_rom[255][15] = 8'd212;
	sample_rom[255][16] = 8'd231;
	sample_rom[255][17] = 8'd231;
	sample_rom[255][18] = 8'd230;
	sample_rom[255][19] = 8'd229;
	sample_rom[255][20] = 8'd228;
	sample_rom[255][21] = 8'd212;
	sample_rom[255][22] = 8'd174;
	sample_rom[255][23] = 8'd162;
	sample_rom[255][24] = 8'd167;
	sample_rom[255][25] = 8'd163;
	sample_rom[255][26] = 8'd146;
	sample_rom[255][27] = 8'd143;
	sample_rom[255][28] = 8'd122;
	sample_rom[255][29] = 8'd80;
	sample_rom[255][30] = 8'd47;
	sample_rom[255][31] = 8'd43;
	sample_rom[255][32] = 8'd67;
	sample_rom[255][33] = 8'd88;
	sample_rom[255][34] = 8'd92;
	sample_rom[255][35] = 8'd101;
	sample_rom[255][36] = 8'd122;
	sample_rom[255][37] = 8'd145;
	sample_rom[255][38] = 8'd157;
	sample_rom[255][39] = 8'd176;
	sample_rom[255][40] = 8'd209;
	sample_rom[255][41] = 8'd225;
	sample_rom[255][42] = 8'd216;
	sample_rom[255][43] = 8'd182;
	sample_rom[255][44] = 8'd162;
	sample_rom[255][45] = 8'd173;
	sample_rom[255][46] = 8'd180;
	sample_rom[255][47] = 8'd161;
	sample_rom[255][48] = 8'd149;
	sample_rom[255][49] = 8'd159;
	sample_rom[255][50] = 8'd164;
	sample_rom[255][51] = 8'd145;
	sample_rom[255][52] = 8'd108;
	sample_rom[255][53] = 8'd87;
	sample_rom[255][54] = 8'd89;
	sample_rom[255][55] = 8'd103;
	sample_rom[255][56] = 8'd101;
	sample_rom[255][57] = 8'd104;
	sample_rom[255][58] = 8'd122;
	sample_rom[255][59] = 8'd99;
	sample_rom[255][60] = 8'd50;
	sample_rom[255][61] = 8'd8;
	sample_rom[255][62] = 8'd1;
	sample_rom[255][63] = 8'd10;
end



endmodule

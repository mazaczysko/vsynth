module bin2bcd (
	input CLK,
	input START,
	input [6:0] bin,
	output reg [8:0] bcd
)



endmodule
